
-- 
-- Definition of  controller
-- 
--      Sun Apr 21 14:19:18 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity controller is
   port (
      clk : IN std_logic ;
      clk_inv : IN std_logic ;
      rst : IN std_logic ;
      initiate : INOUT std_logic ;
      ready_signal : INOUT std_logic ;
      done : INOUT std_logic ;
      enable_mar_in : INOUT std_logic ;
      enable_mdr_in : INOUT std_logic ;
      enable_mdr_out : INOUT std_logic ;
      enable_write : INOUT std_logic ;
      mdr_data_out : INOUT std_logic_vector (255 DOWNTO 0) ;
      label_1_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_2_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_3_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_4_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_5_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_6_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_7_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_8_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_9_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      label_10_output : INOUT std_logic_vector (15 DOWNTO 0) ;
      state : INOUT std_logic_vector (2 DOWNTO 0) ;
      sub_state : INOUT std_logic_vector (2 DOWNTO 0) ;
      answer : OUT std_logic_vector (15 DOWNTO 0) ;
      done_comp : INOUT std_logic) ;
end controller ;

architecture a_controller of controller is
   signal answer_15_EXMPLR, answer_14_EXMPLR, answer_13_EXMPLR, 
      answer_12_EXMPLR, answer_11_EXMPLR, answer_10_EXMPLR, answer_9_EXMPLR, 
      answer_8_EXMPLR, answer_7_EXMPLR, answer_6_EXMPLR, answer_5_EXMPLR, 
      answer_4_EXMPLR, answer_3_EXMPLR, answer_2_EXMPLR, answer_1_EXMPLR, 
      answer_0_EXMPLR, sel_dst_0, nx12877, num_out_2, nx4, nx12879, nx12882, 
      nx12883, nx12885, nx12887, nx20, nx26, nx38, nx56, nx64, 
      enable_decoder_dst_booth, booth_shift_Reg_adder_0_output_17, 
      booth_shift_Reg_adder_0_output_16, booth_shift_Reg_adder_0_output_15, 
      booth_shift_Reg_adder_0_output_14, booth_shift_Reg_adder_0_output_13, 
      booth_shift_Reg_adder_0_output_12, booth_shift_Reg_adder_0_output_11, 
      booth_shift_Reg_adder_0_output_10, booth_shift_Reg_adder_0_output_9, 
      booth_shift_Reg_adder_0_output_8, booth_shift_Reg_adder_0_output_7, 
      booth_shift_Reg_adder_0_output_6, booth_shift_Reg_adder_0_output_5, 
      booth_shift_Reg_adder_0_output_4, booth_shift_Reg_adder_0_output_3, 
      booth_shift_Reg_adder_0_output_2, booth_shift_Reg_adder_0_output_1, 
      booth_shift_Reg_adder_0_output_0, nx12891, nx172, nx12893, nx174, 
      nx186, nx190, nx210, num_in_2, nx242, nx258, nx266, nx278, nx12895, 
      alu_inp1_0, address_out_0, enable_address, nx300, address_in_0, nx320, 
      nx334, nx350, nx358, num_out_0, num_in_0, nx376, nx390, nx412, 
      alu_inp1_1, address_out_1, address_in_1, nx12898, nx414, nx416, 
      num_out_1, num_in_1, nx448, alu_inp1_2, address_out_2, address_in_2, 
      nx464, nx480, nx496, nx516, num_out_3, num_in_3, nx522, alu_inp1_3, 
      address_out_3, address_in_3, nx12901, nx524, nx540, nx548, num_out_4, 
      num_in_4, alu_inp1_4, address_out_4, address_in_4, nx574, nx590, nx606, 
      num_out_5, nx630, alu_inp1_5, address_out_5, address_in_5, nx12905, 
      nx632, nx648, nx656, num_out_6, num_in_6, alu_inp1_6, address_out_6, 
      address_in_6, nx682, nx698, nx714, num_out_7, nx736, alu_inp1_7, 
      address_out_7, address_in_7, nx12907, nx738, nx754, nx12909, nx830, 
      nx846, nx868, nx878, label_4_input_15, label_4_input_state_machine_15, 
      label_4_input_0, booth_booth_integrtaion_3_shift_reg_output_9, 
      booth_booth_integrtaion_3_shift_Reg_count_9, 
      booth_booth_integrtaion_3_shift_Reg_output_8, 
      booth_booth_integrtaion_3_shift_Reg_count_8, 
      booth_booth_integrtaion_3_shift_Reg_output_7, 
      booth_booth_integrtaion_3_shift_Reg_count_7, 
      booth_booth_integrtaion_3_shift_Reg_output_6, 
      booth_booth_integrtaion_3_shift_Reg_count_6, 
      booth_booth_integrtaion_3_shift_Reg_output_5, 
      booth_booth_integrtaion_3_shift_Reg_count_5, 
      booth_booth_integrtaion_3_shift_Reg_output_4, 
      booth_booth_integrtaion_3_shift_Reg_count_4, 
      booth_booth_integrtaion_3_shift_Reg_output_3, 
      booth_booth_integrtaion_3_shift_Reg_count_3, 
      booth_booth_integrtaion_3_shift_Reg_output_2, 
      booth_booth_integrtaion_3_shift_Reg_count_2, 
      booth_booth_integrtaion_3_shift_Reg_output_1, 
      booth_booth_integrtaion_3_shift_Reg_count_1, 
      booth_booth_integrtaion_3_shift_reg_output_0, 
      booth_booth_integrtaion_3_shift_Reg_count_0, 
      booth_booth_integration_output_3_1, booth_booth_integration_output_3_2, 
      booth_booth_integration_output_3_3, booth_booth_integration_output_3_4, 
      booth_booth_integration_output_3_5, booth_booth_integration_output_3_6, 
      booth_booth_integration_output_3_7, booth_booth_integration_output_3_8, 
      booth_booth_integration_output_3_9, 
      booth_booth_integration_output_3_10, 
      booth_booth_integration_output_3_11, 
      booth_booth_integration_output_3_12, 
      booth_booth_integration_output_3_13, 
      booth_booth_integration_output_3_14, 
      booth_booth_integration_output_3_15, 
      booth_booth_integrtaion_3_booth_output_16, nx994, nx1000, 
      booth_booth_integrtaion_3_booth_output_17, nx12913, nx1008, nx1024, 
      booth_booth_integrtaion_3_booth_output_18, nx12915, nx1034, nx1038, 
      nx1052, booth_booth_integrtaion_3_booth_output_19, nx12917, nx1058, 
      nx1062, nx1072, booth_booth_integrtaion_3_booth_output_20, nx12919, 
      nx1082, nx1086, nx1100, booth_booth_integrtaion_3_booth_output_21, 
      nx12921, nx1106, nx1110, nx1120, 
      booth_booth_integrtaion_3_booth_output_22, nx12922, nx1130, nx1134, 
      nx1148, booth_booth_integrtaion_3_booth_output_23, nx12923, nx1154, 
      nx1158, nx1168, booth_booth_integrtaion_3_booth_output_24, nx12925, 
      nx1178, nx1182, nx1196, booth_booth_integrtaion_3_booth_output_25, 
      nx12927, nx1202, nx1206, nx1216, 
      booth_booth_integrtaion_3_booth_output_26, nx12929, nx1226, nx1230, 
      nx1244, booth_booth_integrtaion_3_booth_output_27, nx12930, nx1250, 
      nx1254, nx1264, booth_booth_integrtaion_3_booth_output_28, nx12931, 
      nx1274, nx1278, nx1292, booth_booth_integrtaion_3_booth_output_29, 
      nx12933, nx1298, nx1302, nx1312, 
      booth_booth_integrtaion_3_booth_output_31, nx12935, nx1322, nx1326, 
      nx1340, nx1342, nx1350, nx1356, nx1364, nx1380, nx1388, nx1404, nx1412, 
      nx1428, nx1436, nx1452, nx1460, nx1476, nx1484, nx1500, nx1508, nx1524, 
      nx1530, nx1536, nx1554, nx1566, nx1578, nx1590, nx1602, nx1614, nx1626, 
      nx1638, nx1650, nx1662, nx1674, nx1686, nx1698, nx1710, nx1722, nx1732, 
      label_4_input_state_machine_0, nx1744, label_4_input_1, 
      label_4_input_state_machine_1, nx12939, nx1766, nx1770, 
      label_4_input_2, label_4_input_state_machine_2, nx1798, nx1802, nx1820, 
      label_4_input_3, label_4_input_state_machine_3, nx12943, nx1830, 
      nx1834, label_4_input_4, label_4_input_state_machine_4, nx1862, nx1866, 
      nx1884, label_4_input_5, label_4_input_state_machine_5, nx12946, 
      nx1894, nx1898, label_4_input_6, label_4_input_state_machine_6, nx1926, 
      nx1930, nx1948, label_4_input_7, label_4_input_state_machine_7, 
      nx12949, nx1958, nx1962, label_4_input_8, 
      label_4_input_state_machine_8, nx1990, nx1994, nx2012, label_4_input_9, 
      label_4_input_state_machine_9, nx12953, nx2022, nx2026, 
      label_4_input_10, label_4_input_state_machine_10, nx2054, nx2058, 
      nx2076, label_4_input_11, label_4_input_state_machine_11, nx12955, 
      nx2086, nx2090, label_4_input_12, label_4_input_state_machine_12, 
      nx2118, nx2122, nx2140, label_4_input_13, 
      label_4_input_state_machine_13, nx12959, nx2150, nx2154, 
      label_4_input_14, label_4_input_state_machine_14, nx2182, nx2186, 
      nx2204, nx2208, nx2212, label_3_input_15, 
      label_3_input_state_machine_15, label_3_input_0, 
      booth_booth_integrtaion_2_shift_reg_output_9, 
      booth_booth_integrtaion_2_shift_Reg_count_9, 
      booth_booth_integrtaion_2_shift_Reg_output_8, 
      booth_booth_integrtaion_2_shift_Reg_count_8, 
      booth_booth_integrtaion_2_shift_Reg_output_7, 
      booth_booth_integrtaion_2_shift_Reg_count_7, 
      booth_booth_integrtaion_2_shift_Reg_output_6, 
      booth_booth_integrtaion_2_shift_Reg_count_6, 
      booth_booth_integrtaion_2_shift_Reg_output_5, 
      booth_booth_integrtaion_2_shift_Reg_count_5, 
      booth_booth_integrtaion_2_shift_Reg_output_4, 
      booth_booth_integrtaion_2_shift_Reg_count_4, 
      booth_booth_integrtaion_2_shift_Reg_output_3, 
      booth_booth_integrtaion_2_shift_Reg_count_3, 
      booth_booth_integrtaion_2_shift_Reg_output_2, 
      booth_booth_integrtaion_2_shift_Reg_count_2, 
      booth_booth_integrtaion_2_shift_Reg_output_1, 
      booth_booth_integrtaion_2_shift_Reg_count_1, 
      booth_booth_integrtaion_2_shift_reg_output_0, 
      booth_booth_integrtaion_2_shift_Reg_count_0, 
      booth_booth_integration_output_2_1, booth_booth_integration_output_2_2, 
      booth_booth_integration_output_2_3, booth_booth_integration_output_2_4, 
      booth_booth_integration_output_2_5, booth_booth_integration_output_2_6, 
      booth_booth_integration_output_2_7, booth_booth_integration_output_2_8, 
      booth_booth_integration_output_2_9, 
      booth_booth_integration_output_2_10, 
      booth_booth_integration_output_2_11, 
      booth_booth_integration_output_2_12, 
      booth_booth_integration_output_2_13, 
      booth_booth_integration_output_2_14, 
      booth_booth_integration_output_2_15, 
      booth_booth_integrtaion_2_booth_output_16, nx2332, nx2338, 
      booth_booth_integrtaion_2_booth_output_17, nx12965, nx2346, nx2362, 
      booth_booth_integrtaion_2_booth_output_18, nx12967, nx2372, nx2376, 
      nx2390, booth_booth_integrtaion_2_booth_output_19, nx12969, nx2396, 
      nx2400, nx2410, booth_booth_integrtaion_2_booth_output_20, nx12970, 
      nx2420, nx2424, nx2438, booth_booth_integrtaion_2_booth_output_21, 
      nx12971, nx2444, nx2448, nx2458, 
      booth_booth_integrtaion_2_booth_output_22, nx12973, nx2468, nx2472, 
      nx2486, booth_booth_integrtaion_2_booth_output_23, nx12975, nx2492, 
      nx2496, nx2506, booth_booth_integrtaion_2_booth_output_24, nx12977, 
      nx2516, nx2520, nx2534, booth_booth_integrtaion_2_booth_output_25, 
      nx12978, nx2540, nx2544, nx2554, 
      booth_booth_integrtaion_2_booth_output_26, nx12979, nx2564, nx2568, 
      nx2582, booth_booth_integrtaion_2_booth_output_27, nx12981, nx2588, 
      nx2592, nx2602, booth_booth_integrtaion_2_booth_output_28, nx12983, 
      nx2612, nx2616, nx2630, booth_booth_integrtaion_2_booth_output_29, 
      nx12985, nx2636, nx2640, nx2650, 
      booth_booth_integrtaion_2_booth_output_31, nx12987, nx2660, nx2664, 
      nx2678, nx2680, nx2688, nx2694, nx2702, nx2718, nx2726, nx2742, nx2750, 
      nx2766, nx2774, nx2790, nx2798, nx2814, nx2822, nx2838, nx2846, nx2862, 
      nx2868, nx2874, nx2892, nx2904, nx2916, nx2928, nx2940, nx2952, nx2964, 
      nx2976, nx2988, nx3000, nx3012, nx3024, nx3036, nx3048, nx3060, nx3070, 
      label_3_input_state_machine_0, nx3082, label_3_input_1, 
      label_3_input_state_machine_1, nx12991, nx3104, nx3108, 
      label_3_input_2, label_3_input_state_machine_2, nx3136, nx3140, nx3158, 
      label_3_input_3, label_3_input_state_machine_3, nx12994, nx3168, 
      nx3172, label_3_input_4, label_3_input_state_machine_4, nx3200, nx3204, 
      nx3222, label_3_input_5, label_3_input_state_machine_5, nx12997, 
      nx3232, nx3236, label_3_input_6, label_3_input_state_machine_6, nx3264, 
      nx3268, nx3286, label_3_input_7, label_3_input_state_machine_7, 
      nx13001, nx3296, nx3300, label_3_input_8, 
      label_3_input_state_machine_8, nx3328, nx3332, nx3350, label_3_input_9, 
      label_3_input_state_machine_9, nx13003, nx3360, nx3364, 
      label_3_input_10, label_3_input_state_machine_10, nx3392, nx3396, 
      nx3414, label_3_input_11, label_3_input_state_machine_11, nx13007, 
      nx3424, nx3428, label_3_input_12, label_3_input_state_machine_12, 
      nx3456, nx3460, nx3478, label_3_input_13, 
      label_3_input_state_machine_13, nx13011, nx3488, nx3492, 
      label_3_input_14, label_3_input_state_machine_14, nx3520, nx3524, 
      nx3542, nx3546, nx3550, label_2_input_15, 
      label_2_input_state_machine_15, label_2_input_0, 
      booth_booth_integrtaion_1_shift_reg_output_9, 
      booth_booth_integrtaion_1_shift_Reg_count_9, 
      booth_booth_integrtaion_1_shift_Reg_output_8, 
      booth_booth_integrtaion_1_shift_Reg_count_8, 
      booth_booth_integrtaion_1_shift_Reg_output_7, 
      booth_booth_integrtaion_1_shift_Reg_count_7, 
      booth_booth_integrtaion_1_shift_Reg_output_6, 
      booth_booth_integrtaion_1_shift_Reg_count_6, 
      booth_booth_integrtaion_1_shift_Reg_output_5, 
      booth_booth_integrtaion_1_shift_Reg_count_5, 
      booth_booth_integrtaion_1_shift_Reg_output_4, 
      booth_booth_integrtaion_1_shift_Reg_count_4, 
      booth_booth_integrtaion_1_shift_Reg_output_3, 
      booth_booth_integrtaion_1_shift_Reg_count_3, 
      booth_booth_integrtaion_1_shift_Reg_output_2, 
      booth_booth_integrtaion_1_shift_Reg_count_2, 
      booth_booth_integrtaion_1_shift_Reg_output_1, 
      booth_booth_integrtaion_1_shift_Reg_count_1, 
      booth_booth_integrtaion_1_shift_reg_output_0, 
      booth_booth_integrtaion_1_shift_Reg_count_0, 
      booth_booth_integration_output_1_1, booth_booth_integration_output_1_2, 
      booth_booth_integration_output_1_3, booth_booth_integration_output_1_4, 
      booth_booth_integration_output_1_5, booth_booth_integration_output_1_6, 
      booth_booth_integration_output_1_7, booth_booth_integration_output_1_8, 
      booth_booth_integration_output_1_9, 
      booth_booth_integration_output_1_10, 
      booth_booth_integration_output_1_11, 
      booth_booth_integration_output_1_12, 
      booth_booth_integration_output_1_13, 
      booth_booth_integration_output_1_14, 
      booth_booth_integration_output_1_15, 
      booth_booth_integrtaion_1_booth_output_16, nx3670, nx3676, 
      booth_booth_integrtaion_1_booth_output_17, nx13017, nx3684, nx3700, 
      booth_booth_integrtaion_1_booth_output_18, nx13018, nx3710, nx3714, 
      nx3728, booth_booth_integrtaion_1_booth_output_19, nx13019, nx3734, 
      nx3738, nx3748, booth_booth_integrtaion_1_booth_output_20, nx13021, 
      nx3758, nx3762, nx3776, booth_booth_integrtaion_1_booth_output_21, 
      nx13023, nx3782, nx3786, nx3796, 
      booth_booth_integrtaion_1_booth_output_22, nx13025, nx3806, nx3810, 
      nx3824, booth_booth_integrtaion_1_booth_output_23, nx13026, nx3830, 
      nx3834, nx3844, booth_booth_integrtaion_1_booth_output_24, nx13027, 
      nx3854, nx3858, nx3872, booth_booth_integrtaion_1_booth_output_25, 
      nx13029, nx3878, nx3882, nx3892, 
      booth_booth_integrtaion_1_booth_output_26, nx13031, nx3902, nx3906, 
      nx3920, booth_booth_integrtaion_1_booth_output_27, nx13033, nx3926, 
      nx3930, nx3940, booth_booth_integrtaion_1_booth_output_28, nx13035, 
      nx3950, nx3954, nx3968, booth_booth_integrtaion_1_booth_output_29, 
      nx13037, nx3974, nx3978, nx3988, 
      booth_booth_integrtaion_1_booth_output_31, nx13039, nx3998, nx4002, 
      nx4016, nx4018, nx4026, nx4032, nx4040, nx4056, nx4064, nx4080, nx4088, 
      nx4104, nx4112, nx4128, nx4136, nx4152, nx4160, nx4176, nx4184, nx4200, 
      nx4206, nx4212, nx4230, nx4242, nx4254, nx4266, nx4278, nx4290, nx4302, 
      nx4314, nx4326, nx4338, nx4350, nx4362, nx4374, nx4386, nx4398, nx4408, 
      label_2_input_state_machine_0, nx4420, label_2_input_1, 
      label_2_input_state_machine_1, nx13042, nx4442, nx4446, 
      label_2_input_2, label_2_input_state_machine_2, nx4474, nx4478, nx4496, 
      label_2_input_3, label_2_input_state_machine_3, nx13045, nx4506, 
      nx4510, label_2_input_4, label_2_input_state_machine_4, nx4538, nx4542, 
      nx4560, label_2_input_5, label_2_input_state_machine_5, nx13049, 
      nx4570, nx4574, label_2_input_6, label_2_input_state_machine_6, nx4602, 
      nx4606, nx4624, label_2_input_7, label_2_input_state_machine_7, 
      nx13051, nx4634, nx4638, label_2_input_8, 
      label_2_input_state_machine_8, nx4666, nx4670, nx4688, label_2_input_9, 
      label_2_input_state_machine_9, nx13055, nx4698, nx4702, 
      label_2_input_10, label_2_input_state_machine_10, nx4730, nx4734, 
      nx4752, label_2_input_11, label_2_input_state_machine_11, nx13059, 
      nx4762, nx4766, label_2_input_12, label_2_input_state_machine_12, 
      nx4794, nx4798, nx4816, label_2_input_13, 
      label_2_input_state_machine_13, nx13063, nx4826, nx4830, 
      label_2_input_14, label_2_input_state_machine_14, nx4858, nx4862, 
      nx4880, nx4884, nx4888, label_1_input_15, 
      label_1_input_state_machine_15, label_1_input_0, 
      booth_booth_integrtaion_0_shift_reg_output_9, 
      booth_booth_integrtaion_0_shift_Reg_count_9, 
      booth_booth_integrtaion_0_shift_Reg_output_8, 
      booth_booth_integrtaion_0_shift_Reg_count_8, 
      booth_booth_integrtaion_0_shift_Reg_output_7, 
      booth_booth_integrtaion_0_shift_Reg_count_7, 
      booth_booth_integrtaion_0_shift_Reg_output_6, 
      booth_booth_integrtaion_0_shift_Reg_count_6, 
      booth_booth_integrtaion_0_shift_Reg_output_5, 
      booth_booth_integrtaion_0_shift_Reg_count_5, 
      booth_booth_integrtaion_0_shift_Reg_output_4, 
      booth_booth_integrtaion_0_shift_Reg_count_4, 
      booth_booth_integrtaion_0_shift_Reg_output_3, 
      booth_booth_integrtaion_0_shift_Reg_count_3, 
      booth_booth_integrtaion_0_shift_Reg_output_2, 
      booth_booth_integrtaion_0_shift_Reg_count_2, 
      booth_booth_integrtaion_0_shift_Reg_output_1, 
      booth_booth_integrtaion_0_shift_Reg_count_1, 
      booth_booth_integrtaion_0_shift_reg_output_0, 
      booth_booth_integrtaion_0_shift_Reg_count_0, 
      booth_booth_integration_output_0_1, booth_booth_integration_output_0_2, 
      booth_booth_integration_output_0_3, booth_booth_integration_output_0_4, 
      booth_booth_integration_output_0_5, booth_booth_integration_output_0_6, 
      booth_booth_integration_output_0_7, booth_booth_integration_output_0_8, 
      booth_booth_integration_output_0_9, 
      booth_booth_integration_output_0_10, 
      booth_booth_integration_output_0_11, 
      booth_booth_integration_output_0_12, 
      booth_booth_integration_output_0_13, 
      booth_booth_integration_output_0_14, 
      booth_booth_integration_output_0_15, 
      booth_booth_integrtaion_0_booth_output_16, nx5008, nx5014, 
      booth_booth_integrtaion_0_booth_output_17, nx13067, nx5022, nx5038, 
      booth_booth_integrtaion_0_booth_output_18, nx13069, nx5048, nx5052, 
      nx5066, booth_booth_integrtaion_0_booth_output_19, nx13071, nx5072, 
      nx5076, nx5086, booth_booth_integrtaion_0_booth_output_20, nx13073, 
      nx5096, nx5100, nx5114, booth_booth_integrtaion_0_booth_output_21, 
      nx13074, nx5120, nx5124, nx5134, 
      booth_booth_integrtaion_0_booth_output_22, nx13075, nx5144, nx5148, 
      nx5162, booth_booth_integrtaion_0_booth_output_23, nx13077, nx5168, 
      nx5172, nx5182, booth_booth_integrtaion_0_booth_output_24, nx13079, 
      nx5192, nx5196, nx5210, booth_booth_integrtaion_0_booth_output_25, 
      nx13081, nx5216, nx5220, nx5230, 
      booth_booth_integrtaion_0_booth_output_26, nx13083, nx5240, nx5244, 
      nx5258, booth_booth_integrtaion_0_booth_output_27, nx13085, nx5264, 
      nx5268, nx5278, booth_booth_integrtaion_0_booth_output_28, nx13087, 
      nx5288, nx5292, nx5306, booth_booth_integrtaion_0_booth_output_29, 
      nx13089, nx5312, nx5316, nx5326, 
      booth_booth_integrtaion_0_booth_output_31, nx13090, nx5336, nx5340, 
      nx5354, nx5356, nx5364, nx5370, nx5378, nx5394, nx5402, nx5418, nx5426, 
      nx5442, nx5450, nx5466, nx5474, nx5490, nx5498, nx5514, nx5522, nx5538, 
      nx5544, nx5550, nx5568, nx5580, nx5592, nx5604, nx5616, nx5628, nx5640, 
      nx5652, nx5664, nx5676, nx5688, nx5700, nx5712, nx5724, nx5736, nx5746, 
      label_1_input_state_machine_0, nx5758, label_1_input_1, 
      label_1_input_state_machine_1, nx13093, nx5780, nx5784, 
      label_1_input_2, label_1_input_state_machine_2, nx5812, nx5816, nx5834, 
      label_1_input_3, label_1_input_state_machine_3, nx13097, nx5844, 
      nx5848, label_1_input_4, label_1_input_state_machine_4, nx5876, nx5880, 
      nx5898, label_1_input_5, label_1_input_state_machine_5, nx13099, 
      nx5908, nx5912, label_1_input_6, label_1_input_state_machine_6, nx5940, 
      nx5944, nx5962, label_1_input_7, label_1_input_state_machine_7, 
      nx13103, nx5972, nx5976, label_1_input_8, 
      label_1_input_state_machine_8, nx6004, nx6008, nx6026, label_1_input_9, 
      label_1_input_state_machine_9, nx13107, nx6036, nx6040, 
      label_1_input_10, label_1_input_state_machine_10, nx6068, nx6072, 
      nx6090, label_1_input_11, label_1_input_state_machine_11, nx13111, 
      nx6100, nx6104, label_1_input_12, label_1_input_state_machine_12, 
      nx6132, nx6136, nx6154, label_1_input_13, 
      label_1_input_state_machine_13, nx13114, nx6164, nx6168, 
      label_1_input_14, label_1_input_state_machine_14, nx6196, nx6200, 
      nx6218, nx6222, nx6226, max_calc_state_2, max_calc_start, start_comp, 
      nx6244, max_calc_state_0, max_calc_state_3, max_calc_state_1, nx6300, 
      nx6342, max_calc_comparator_first_inp1_0, nx6352, max_calc_ans1_0, 
      nx6368, nx13121, nx6388, max_calc_ans6_0, max_calc_ans5_0, 
      max_calc_comparator_fifth_inp1_0, label_9_input_0, 
      booth_booth_integrtaion_8_shift_reg_output_9, 
      booth_booth_integrtaion_8_shift_Reg_count_9, 
      booth_booth_integrtaion_8_shift_Reg_output_8, 
      booth_booth_integrtaion_8_shift_Reg_count_8, 
      booth_booth_integrtaion_8_shift_Reg_output_7, 
      booth_booth_integrtaion_8_shift_Reg_count_7, 
      booth_booth_integrtaion_8_shift_Reg_output_6, 
      booth_booth_integrtaion_8_shift_Reg_count_6, 
      booth_booth_integrtaion_8_shift_Reg_output_5, 
      booth_booth_integrtaion_8_shift_Reg_count_5, 
      booth_booth_integrtaion_8_shift_Reg_output_4, 
      booth_booth_integrtaion_8_shift_Reg_count_4, 
      booth_booth_integrtaion_8_shift_Reg_output_3, 
      booth_booth_integrtaion_8_shift_Reg_count_3, 
      booth_booth_integrtaion_8_shift_Reg_output_2, 
      booth_booth_integrtaion_8_shift_Reg_count_2, 
      booth_booth_integrtaion_8_shift_Reg_output_1, 
      booth_booth_integrtaion_8_shift_Reg_count_1, 
      booth_booth_integrtaion_8_shift_reg_output_0, 
      booth_booth_integrtaion_8_shift_Reg_count_0, 
      booth_booth_integration_output_8_1, booth_booth_integration_output_8_2, 
      booth_booth_integration_output_8_3, booth_booth_integration_output_8_4, 
      booth_booth_integration_output_8_5, booth_booth_integration_output_8_6, 
      booth_booth_integration_output_8_7, booth_booth_integration_output_8_8, 
      booth_booth_integration_output_8_9, 
      booth_booth_integration_output_8_10, 
      booth_booth_integration_output_8_11, 
      booth_booth_integration_output_8_12, 
      booth_booth_integration_output_8_13, 
      booth_booth_integration_output_8_14, 
      booth_booth_integration_output_8_15, 
      booth_booth_integrtaion_8_booth_output_16, nx6508, nx6514, 
      booth_booth_integrtaion_8_booth_output_17, nx13123, nx6522, nx6538, 
      booth_booth_integrtaion_8_booth_output_18, nx13125, nx6548, nx6552, 
      nx6566, booth_booth_integrtaion_8_booth_output_19, nx13127, nx6572, 
      nx6576, nx6586, booth_booth_integrtaion_8_booth_output_20, nx13129, 
      nx6596, nx6600, nx6614, booth_booth_integrtaion_8_booth_output_21, 
      nx13131, nx6620, nx6624, nx6634, 
      booth_booth_integrtaion_8_booth_output_22, nx13133, nx6644, nx6648, 
      nx6662, booth_booth_integrtaion_8_booth_output_23, nx13135, nx6668, 
      nx6672, nx6682, booth_booth_integrtaion_8_booth_output_24, nx13137, 
      nx6692, nx6696, nx6710, booth_booth_integrtaion_8_booth_output_25, 
      nx13138, nx6716, nx6720, nx6730, 
      booth_booth_integrtaion_8_booth_output_26, nx13139, nx6740, nx6744, 
      nx6758, booth_booth_integrtaion_8_booth_output_27, nx13141, nx6764, 
      nx6768, nx6778, booth_booth_integrtaion_8_booth_output_28, nx13143, 
      nx6788, nx6792, nx6806, booth_booth_integrtaion_8_booth_output_29, 
      nx13145, nx6812, nx6816, nx6826, 
      booth_booth_integrtaion_8_booth_output_31, nx13146, nx6836, nx6840, 
      nx6854, nx6856, nx6864, nx6870, nx6878, nx6894, nx6902, nx6918, nx6926, 
      nx6942, nx6950, nx6966, nx6974, nx6990, nx6998, nx7014, nx7022, nx7038, 
      nx7044, nx7050, nx7068, nx7080, nx7092, nx7104, nx7116, nx7128, nx7140, 
      nx7152, nx7164, nx7176, nx7188, nx7200, nx7212, nx7224, nx7236, nx7248, 
      label_9_input_state_machine_0, nx7260, label_10_input_14, 
      label_10_input_state_machine_14, label_10_input_0, 
      booth_booth_integrtaion_9_shift_reg_output_9, 
      booth_booth_integrtaion_9_shift_Reg_count_9, 
      booth_booth_integrtaion_9_shift_Reg_output_8, 
      booth_booth_integrtaion_9_shift_Reg_count_8, 
      booth_booth_integrtaion_9_shift_Reg_output_7, 
      booth_booth_integrtaion_9_shift_Reg_count_7, 
      booth_booth_integrtaion_9_shift_Reg_output_6, 
      booth_booth_integrtaion_9_shift_Reg_count_6, 
      booth_booth_integrtaion_9_shift_Reg_output_5, 
      booth_booth_integrtaion_9_shift_Reg_count_5, 
      booth_booth_integrtaion_9_shift_Reg_output_4, 
      booth_booth_integrtaion_9_shift_Reg_count_4, 
      booth_booth_integrtaion_9_shift_Reg_output_3, 
      booth_booth_integrtaion_9_shift_Reg_count_3, 
      booth_booth_integrtaion_9_shift_Reg_output_2, 
      booth_booth_integrtaion_9_shift_Reg_count_2, 
      booth_booth_integrtaion_9_shift_Reg_output_1, 
      booth_booth_integrtaion_9_shift_Reg_count_1, 
      booth_booth_integrtaion_9_shift_reg_output_0, 
      booth_booth_integrtaion_9_shift_Reg_count_0, 
      booth_booth_integration_output_9_1, booth_booth_integration_output_9_2, 
      booth_booth_integration_output_9_3, booth_booth_integration_output_9_4, 
      booth_booth_integration_output_9_5, booth_booth_integration_output_9_6, 
      booth_booth_integration_output_9_7, booth_booth_integration_output_9_8, 
      booth_booth_integration_output_9_9, 
      booth_booth_integration_output_9_10, 
      booth_booth_integration_output_9_11, 
      booth_booth_integration_output_9_12, 
      booth_booth_integration_output_9_13, 
      booth_booth_integration_output_9_14, 
      booth_booth_integration_output_9_15, 
      booth_booth_integrtaion_9_booth_output_16, nx7388, nx7394, 
      booth_booth_integrtaion_9_booth_output_17, nx13149, nx7402, nx7418, 
      booth_booth_integrtaion_9_booth_output_18, nx13151, nx7428, nx7432, 
      nx7446, booth_booth_integrtaion_9_booth_output_19, nx13153, nx7452, 
      nx7456, nx7466, booth_booth_integrtaion_9_booth_output_20, nx13155, 
      nx7476, nx7480, nx7494, booth_booth_integrtaion_9_booth_output_21, 
      nx13157, nx7500, nx7504, nx7514, 
      booth_booth_integrtaion_9_booth_output_22, nx13159, nx7524, nx7528, 
      nx7542, booth_booth_integrtaion_9_booth_output_23, nx13161, nx7548, 
      nx7552, nx7562, booth_booth_integrtaion_9_booth_output_24, nx13162, 
      nx7572, nx7576, nx7590, booth_booth_integrtaion_9_booth_output_25, 
      nx13163, nx7596, nx7600, nx7610, 
      booth_booth_integrtaion_9_booth_output_26, nx13165, nx7620, nx7624, 
      nx7638, booth_booth_integrtaion_9_booth_output_27, nx13167, nx7644, 
      nx7648, nx7658, booth_booth_integrtaion_9_booth_output_28, nx13169, 
      nx7668, nx7672, nx7686, booth_booth_integrtaion_9_booth_output_29, 
      nx13170, nx7692, nx7696, nx7706, 
      booth_booth_integrtaion_9_booth_output_31, nx13171, nx7716, nx7720, 
      nx7734, nx7736, nx7744, nx7750, nx7758, nx7774, nx7782, nx7798, nx7806, 
      nx7822, nx7830, nx7846, nx7854, nx7870, nx7878, nx7894, nx7902, nx7918, 
      nx7924, nx7930, nx7948, nx7960, nx7972, nx7984, nx7996, nx8008, nx8020, 
      nx8032, nx8044, nx8056, nx8068, nx8080, nx8092, nx8104, nx8116, nx8126, 
      label_10_input_state_machine_0, nx8138, label_10_input_1, 
      label_10_input_state_machine_1, nx13175, nx8160, nx8164, 
      label_10_input_2, label_10_input_state_machine_2, nx8192, nx8196, 
      nx8214, label_10_input_3, label_10_input_state_machine_3, nx13179, 
      nx8224, nx8228, label_10_input_4, label_10_input_state_machine_4, 
      nx8256, nx8260, nx8278, label_10_input_5, 
      label_10_input_state_machine_5, nx13183, nx8288, nx8292, 
      label_10_input_6, label_10_input_state_machine_6, nx8320, nx8324, 
      nx8342, label_10_input_7, label_10_input_state_machine_7, nx13187, 
      nx8352, nx8356, label_10_input_8, label_10_input_state_machine_8, 
      nx8384, nx8388, nx8406, label_10_input_9, 
      label_10_input_state_machine_9, nx13191, nx8416, nx8420, 
      label_10_input_10, label_10_input_state_machine_10, nx8448, nx8452, 
      nx8470, label_10_input_11, label_10_input_state_machine_11, nx13195, 
      nx8480, nx8484, label_10_input_12, label_10_input_state_machine_12, 
      nx8512, nx8516, nx8534, label_10_input_13, 
      label_10_input_state_machine_13, nx13199, nx8544, nx8548, nx8570, 
      nx8574, max_calc_comparator_fifth_inp1_14, label_9_input_14, 
      label_9_input_state_machine_14, label_9_input_1, 
      label_9_input_state_machine_1, nx13200, nx8610, nx8614, 
      label_9_input_2, label_9_input_state_machine_2, nx8642, nx8646, nx8664, 
      label_9_input_3, label_9_input_state_machine_3, nx13202, nx8674, 
      nx8678, label_9_input_4, label_9_input_state_machine_4, nx8706, nx8710, 
      nx8728, label_9_input_5, label_9_input_state_machine_5, nx13204, 
      nx8738, nx8742, label_9_input_6, label_9_input_state_machine_6, nx8770, 
      nx8774, nx8792, label_9_input_7, label_9_input_state_machine_7, 
      nx13207, nx8802, nx8806, label_9_input_8, 
      label_9_input_state_machine_8, nx8834, nx8838, nx8856, label_9_input_9, 
      label_9_input_state_machine_9, nx13211, nx8866, nx8870, 
      label_9_input_10, label_9_input_state_machine_10, nx8898, nx8902, 
      nx8920, label_9_input_11, label_9_input_state_machine_11, nx13213, 
      nx8930, nx8934, label_9_input_12, label_9_input_state_machine_12, 
      nx8962, nx8966, nx8984, label_9_input_13, 
      label_9_input_state_machine_13, nx13215, nx8994, nx8998, nx9020, 
      nx9024, nx9044, max_calc_comparator_fifth_inp2_13, 
      max_calc_comparator_fifth_inp1_13, max_calc_comparator_fifth_inp1_12, 
      nx9080, max_calc_comparator_fifth_inp2_11, 
      max_calc_comparator_fifth_inp1_11, max_calc_comparator_fifth_inp1_10, 
      nx9116, max_calc_comparator_fifth_inp2_9, 
      max_calc_comparator_fifth_inp1_9, max_calc_comparator_fifth_inp1_8, 
      nx9152, max_calc_comparator_fifth_inp2_7, 
      max_calc_comparator_fifth_inp1_7, max_calc_comparator_fifth_inp1_6, 
      nx9188, max_calc_comparator_fifth_inp2_5, 
      max_calc_comparator_fifth_inp1_5, max_calc_comparator_fifth_inp1_4, 
      nx9224, max_calc_comparator_fifth_inp2_3, 
      max_calc_comparator_fifth_inp1_3, max_calc_comparator_fifth_inp1_2, 
      nx9260, max_calc_comparator_fifth_inp2_1, nx9278, nx9302, nx9318, 
      nx9334, nx9350, nx9366, nx9382, nx9398, label_10_input_15, 
      label_10_input_state_machine_15, nx9420, nx9424, nx9428, 
      label_9_input_15, label_9_input_state_machine_15, nx9460, nx9464, 
      nx9468, nx9488, nx9490, nx9498, nx9508, nx9512, 
      max_calc_comparator_first_inp2_14, max_calc_ans2_14, 
      max_calc_comparator_second_inp1_14, max_calc_ans3_14, 
      max_calc_comparator_third_inp1_14, label_5_input_14, 
      label_5_input_state_machine_14, label_5_input_0, 
      booth_booth_integrtaion_4_shift_reg_output_9, 
      booth_booth_integrtaion_4_shift_Reg_count_9, 
      booth_booth_integrtaion_4_shift_Reg_output_8, 
      booth_booth_integrtaion_4_shift_Reg_count_8, 
      booth_booth_integrtaion_4_shift_Reg_output_7, 
      booth_booth_integrtaion_4_shift_Reg_count_7, 
      booth_booth_integrtaion_4_shift_Reg_output_6, 
      booth_booth_integrtaion_4_shift_Reg_count_6, 
      booth_booth_integrtaion_4_shift_Reg_output_5, 
      booth_booth_integrtaion_4_shift_Reg_count_5, 
      booth_booth_integrtaion_4_shift_Reg_output_4, 
      booth_booth_integrtaion_4_shift_Reg_count_4, 
      booth_booth_integrtaion_4_shift_Reg_output_3, 
      booth_booth_integrtaion_4_shift_Reg_count_3, 
      booth_booth_integrtaion_4_shift_Reg_output_2, 
      booth_booth_integrtaion_4_shift_Reg_count_2, 
      booth_booth_integrtaion_4_shift_Reg_output_1, 
      booth_booth_integrtaion_4_shift_Reg_count_1, 
      booth_booth_integrtaion_4_shift_reg_output_0, 
      booth_booth_integrtaion_4_shift_Reg_count_0, 
      booth_booth_integration_output_4_1, booth_booth_integration_output_4_2, 
      booth_booth_integration_output_4_3, booth_booth_integration_output_4_4, 
      booth_booth_integration_output_4_5, booth_booth_integration_output_4_6, 
      booth_booth_integration_output_4_7, booth_booth_integration_output_4_8, 
      booth_booth_integration_output_4_9, 
      booth_booth_integration_output_4_10, 
      booth_booth_integration_output_4_11, 
      booth_booth_integration_output_4_12, 
      booth_booth_integration_output_4_13, 
      booth_booth_integration_output_4_14, 
      booth_booth_integration_output_4_15, 
      booth_booth_integrtaion_4_booth_output_16, nx9646, nx9652, 
      booth_booth_integrtaion_4_booth_output_17, nx13217, nx9660, nx9676, 
      booth_booth_integrtaion_4_booth_output_18, nx13219, nx9686, nx9690, 
      nx9704, booth_booth_integrtaion_4_booth_output_19, nx13221, nx9710, 
      nx9714, nx9724, booth_booth_integrtaion_4_booth_output_20, nx13223, 
      nx9734, nx9738, nx9752, booth_booth_integrtaion_4_booth_output_21, 
      nx13224, nx9758, nx9762, nx9772, 
      booth_booth_integrtaion_4_booth_output_22, nx13225, nx9782, nx9786, 
      nx9800, booth_booth_integrtaion_4_booth_output_23, nx13226, nx9806, 
      nx9810, nx9820, booth_booth_integrtaion_4_booth_output_24, nx13227, 
      nx9830, nx9834, nx9848, booth_booth_integrtaion_4_booth_output_25, 
      nx13228, nx9854, nx9858, nx9868, 
      booth_booth_integrtaion_4_booth_output_26, nx13229, nx9878, nx9882, 
      nx9896, booth_booth_integrtaion_4_booth_output_27, nx13231, nx9902, 
      nx9906, nx9916, booth_booth_integrtaion_4_booth_output_28, nx13233, 
      nx9926, nx9930, nx9944, booth_booth_integrtaion_4_booth_output_29, 
      nx13235, nx9950, nx9954, nx9964, 
      booth_booth_integrtaion_4_booth_output_31, nx13236, nx9974, nx9978, 
      nx9992, nx9994, nx10002, nx10008, nx10016, nx10032, nx10040, nx10056, 
      nx10064, nx10080, nx10088, nx10104, nx10112, nx10128, nx10136, nx10152, 
      nx10160, nx10176, nx10182, nx10188, nx10206, nx10218, nx10230, nx10242, 
      nx10254, nx10266, nx10278, nx10290, nx10302, nx10314, nx10326, nx10338, 
      nx10350, nx10362, nx10374, nx10384, label_5_input_state_machine_0, 
      nx10396, label_5_input_1, label_5_input_state_machine_1, nx13238, 
      nx10418, nx10422, label_5_input_2, label_5_input_state_machine_2, 
      nx10450, nx10454, nx10472, label_5_input_3, 
      label_5_input_state_machine_3, nx13240, nx10482, nx10486, 
      label_5_input_4, label_5_input_state_machine_4, nx10514, nx10518, 
      nx10536, label_5_input_5, label_5_input_state_machine_5, nx13243, 
      nx10546, nx10550, label_5_input_6, label_5_input_state_machine_6, 
      nx10578, nx10582, nx10600, label_5_input_7, 
      label_5_input_state_machine_7, nx13247, nx10610, nx10614, 
      label_5_input_8, label_5_input_state_machine_8, nx10642, nx10646, 
      nx10664, label_5_input_9, label_5_input_state_machine_9, nx13249, 
      nx10674, nx10678, label_5_input_10, label_5_input_state_machine_10, 
      nx10706, nx10710, nx10728, label_5_input_11, 
      label_5_input_state_machine_11, nx13251, nx10738, nx10742, 
      label_5_input_12, label_5_input_state_machine_12, nx10770, nx10774, 
      nx10792, label_5_input_13, label_5_input_state_machine_13, nx13253, 
      nx10802, nx10806, nx10828, nx10832, label_6_input_14, 
      label_6_input_state_machine_14, label_6_input_0, 
      booth_booth_integrtaion_5_shift_reg_output_9, 
      booth_booth_integrtaion_5_shift_Reg_count_9, 
      booth_booth_integrtaion_5_shift_Reg_output_8, 
      booth_booth_integrtaion_5_shift_Reg_count_8, 
      booth_booth_integrtaion_5_shift_Reg_output_7, 
      booth_booth_integrtaion_5_shift_Reg_count_7, 
      booth_booth_integrtaion_5_shift_Reg_output_6, 
      booth_booth_integrtaion_5_shift_Reg_count_6, 
      booth_booth_integrtaion_5_shift_Reg_output_5, 
      booth_booth_integrtaion_5_shift_Reg_count_5, 
      booth_booth_integrtaion_5_shift_Reg_output_4, 
      booth_booth_integrtaion_5_shift_Reg_count_4, 
      booth_booth_integrtaion_5_shift_Reg_output_3, 
      booth_booth_integrtaion_5_shift_Reg_count_3, 
      booth_booth_integrtaion_5_shift_Reg_output_2, 
      booth_booth_integrtaion_5_shift_Reg_count_2, 
      booth_booth_integrtaion_5_shift_Reg_output_1, 
      booth_booth_integrtaion_5_shift_Reg_count_1, 
      booth_booth_integrtaion_5_shift_reg_output_0, 
      booth_booth_integrtaion_5_shift_Reg_count_0, 
      booth_booth_integration_output_5_1, booth_booth_integration_output_5_2, 
      booth_booth_integration_output_5_3, booth_booth_integration_output_5_4, 
      booth_booth_integration_output_5_5, booth_booth_integration_output_5_6, 
      booth_booth_integration_output_5_7, booth_booth_integration_output_5_8, 
      booth_booth_integration_output_5_9, 
      booth_booth_integration_output_5_10, 
      booth_booth_integration_output_5_11, 
      booth_booth_integration_output_5_12, 
      booth_booth_integration_output_5_13, 
      booth_booth_integration_output_5_14, 
      booth_booth_integration_output_5_15, 
      booth_booth_integrtaion_5_booth_output_16, nx10968, nx10974, 
      booth_booth_integrtaion_5_booth_output_17, nx13257, nx10982, nx10998, 
      booth_booth_integrtaion_5_booth_output_18, nx13259, nx11008, nx11012, 
      nx11026, booth_booth_integrtaion_5_booth_output_19, nx13260, nx11032, 
      nx11036, nx11046, booth_booth_integrtaion_5_booth_output_20, nx13261, 
      nx11056, nx11060, nx11074, booth_booth_integrtaion_5_booth_output_21, 
      nx13262, nx11080, nx11084, nx11094, 
      booth_booth_integrtaion_5_booth_output_22, nx13263, nx11104, nx11108, 
      nx11122, booth_booth_integrtaion_5_booth_output_23, nx13264, nx11128, 
      nx11132, nx11142, booth_booth_integrtaion_5_booth_output_24, nx13265, 
      nx11152, nx11156, nx11170, booth_booth_integrtaion_5_booth_output_25, 
      nx13267, nx11176, nx11180, nx11190, 
      booth_booth_integrtaion_5_booth_output_26, nx13269, nx11200, nx11204, 
      nx11218, booth_booth_integrtaion_5_booth_output_27, nx13271, nx11224, 
      nx11228, nx11238, booth_booth_integrtaion_5_booth_output_28, nx13272, 
      nx11248, nx11252, nx11266, booth_booth_integrtaion_5_booth_output_29, 
      nx13273, nx11272, nx11276, nx11286, 
      booth_booth_integrtaion_5_booth_output_31, nx13274, nx11296, nx11300, 
      nx11314, nx11316, nx11324, nx11330, nx11338, nx11354, nx11362, nx11378, 
      nx11386, nx11402, nx11410, nx11426, nx11434, nx11450, nx11458, nx11474, 
      nx11482, nx11498, nx11504, nx11510, nx11528, nx11540, nx11552, nx11564, 
      nx11576, nx11588, nx11600, nx11612, nx11624, nx11636, nx11648, nx11660, 
      nx11672, nx11684, nx11696, nx11706, label_6_input_state_machine_0, 
      nx11718, label_6_input_1, label_6_input_state_machine_1, nx13276, 
      nx11740, nx11744, label_6_input_2, label_6_input_state_machine_2, 
      nx11772, nx11776, nx11794, label_6_input_3, 
      label_6_input_state_machine_3, nx13279, nx11804, nx11808, 
      label_6_input_4, label_6_input_state_machine_4, nx11836, nx11840, 
      nx11858, label_6_input_5, label_6_input_state_machine_5, nx13283, 
      nx11868, nx11872, label_6_input_6, label_6_input_state_machine_6, 
      nx11900, nx11904, nx11922, label_6_input_7, 
      label_6_input_state_machine_7, nx13285, nx11932, nx11936, 
      label_6_input_8, label_6_input_state_machine_8, nx11964, nx11968, 
      nx11986, label_6_input_9, label_6_input_state_machine_9, nx13287, 
      nx11996, nx12000, label_6_input_10, label_6_input_state_machine_10, 
      nx12028, nx12032, nx12050, label_6_input_11, 
      label_6_input_state_machine_11, nx13289, nx12060, nx12064, 
      label_6_input_12, label_6_input_state_machine_12, nx12092, nx12096, 
      nx12114, label_6_input_13, label_6_input_state_machine_13, nx13293, 
      nx12124, nx12128, nx12150, nx12154, nx12176, 
      max_calc_comparator_third_inp2_13, max_calc_comparator_third_inp1_13, 
      max_calc_comparator_third_inp1_12, nx12220, 
      max_calc_comparator_third_inp2_11, max_calc_comparator_third_inp1_11, 
      max_calc_comparator_third_inp1_10, nx12264, 
      max_calc_comparator_third_inp2_9, max_calc_comparator_third_inp1_9, 
      max_calc_comparator_third_inp1_8, nx12308, 
      max_calc_comparator_third_inp2_7, max_calc_comparator_third_inp1_7, 
      max_calc_comparator_third_inp1_6, nx12352, 
      max_calc_comparator_third_inp2_5, max_calc_comparator_third_inp1_5, 
      max_calc_comparator_third_inp1_4, nx12396, 
      max_calc_comparator_third_inp2_3, max_calc_comparator_third_inp1_3, 
      max_calc_comparator_third_inp1_2, nx12440, 
      max_calc_comparator_third_inp2_1, nx12462, 
      max_calc_comparator_third_inp1_0, nx12498, nx12514, nx12530, nx12546, 
      nx12562, nx12578, nx12594, label_6_input_15, 
      label_6_input_state_machine_15, nx12616, nx12620, nx12624, 
      label_5_input_15, label_5_input_state_machine_15, nx12658, nx12662, 
      nx12666, nx12688, nx12690, nx12712, max_calc_ans4_14, 
      max_calc_comparator_fourth_inp1_14, label_7_input_14, 
      label_7_input_state_machine_14, label_7_input_0, 
      booth_booth_integrtaion_6_shift_reg_output_9, 
      booth_booth_integrtaion_6_shift_Reg_count_9, 
      booth_booth_integrtaion_6_shift_Reg_output_8, 
      booth_booth_integrtaion_6_shift_Reg_count_8, 
      booth_booth_integrtaion_6_shift_Reg_output_7, 
      booth_booth_integrtaion_6_shift_Reg_count_7, 
      booth_booth_integrtaion_6_shift_Reg_output_6, 
      booth_booth_integrtaion_6_shift_Reg_count_6, 
      booth_booth_integrtaion_6_shift_Reg_output_5, 
      booth_booth_integrtaion_6_shift_Reg_count_5, 
      booth_booth_integrtaion_6_shift_Reg_output_4, 
      booth_booth_integrtaion_6_shift_Reg_count_4, 
      booth_booth_integrtaion_6_shift_Reg_output_3, 
      booth_booth_integrtaion_6_shift_Reg_count_3, 
      booth_booth_integrtaion_6_shift_Reg_output_2, 
      booth_booth_integrtaion_6_shift_Reg_count_2, 
      booth_booth_integrtaion_6_shift_Reg_output_1, 
      booth_booth_integrtaion_6_shift_Reg_count_1, 
      booth_booth_integrtaion_6_shift_reg_output_0, 
      booth_booth_integrtaion_6_shift_Reg_count_0, 
      booth_booth_integration_output_6_1, booth_booth_integration_output_6_2, 
      booth_booth_integration_output_6_3, booth_booth_integration_output_6_4, 
      booth_booth_integration_output_6_5, booth_booth_integration_output_6_6, 
      booth_booth_integration_output_6_7, booth_booth_integration_output_6_8, 
      booth_booth_integration_output_6_9, 
      booth_booth_integration_output_6_10, 
      booth_booth_integration_output_6_11, 
      booth_booth_integration_output_6_12, 
      booth_booth_integration_output_6_13, 
      booth_booth_integration_output_6_14, 
      booth_booth_integration_output_6_15, 
      booth_booth_integrtaion_6_booth_output_16, nx12836, nx12842, 
      booth_booth_integrtaion_6_booth_output_17, nx13296, nx12850, nx12866, 
      booth_booth_integrtaion_6_booth_output_18, nx13297, nx12876, nx12880, 
      nx12894, booth_booth_integrtaion_6_booth_output_19, nx13298, nx12900, 
      nx12904, nx12914, booth_booth_integrtaion_6_booth_output_20, nx13299, 
      nx12924, nx12928, nx12942, booth_booth_integrtaion_6_booth_output_21, 
      nx13300, nx12948, nx12952, nx12962, 
      booth_booth_integrtaion_6_booth_output_22, nx13301, nx12972, nx12976, 
      nx12990, booth_booth_integrtaion_6_booth_output_23, nx13303, nx12996, 
      nx13000, nx13010, booth_booth_integrtaion_6_booth_output_24, nx13305, 
      nx13020, nx13024, nx13038, booth_booth_integrtaion_6_booth_output_25, 
      nx13307, nx13044, nx13048, nx13058, 
      booth_booth_integrtaion_6_booth_output_26, nx13308, nx13068, nx13072, 
      nx13086, booth_booth_integrtaion_6_booth_output_27, nx13309, nx13092, 
      nx13096, nx13106, booth_booth_integrtaion_6_booth_output_28, nx13310, 
      nx13116, nx13120, nx13134, booth_booth_integrtaion_6_booth_output_29, 
      nx13311, nx13140, nx13144, nx13154, 
      booth_booth_integrtaion_6_booth_output_31, nx13312, nx13164, nx13168, 
      nx13182, nx13184, nx13192, nx13198, nx13206, nx13222, nx13230, nx13246, 
      nx13254, nx13270, nx13278, nx13294, nx13302, nx13318, nx13326, nx13342, 
      nx13350, nx13366, nx13372, nx13378, nx13396, nx13408, nx13420, nx13432, 
      nx13444, nx13456, nx13468, nx13480, nx13492, nx13504, nx13516, nx13528, 
      nx13540, nx13552, nx13564, nx13574, label_7_input_state_machine_0, 
      nx13586, label_7_input_1, label_7_input_state_machine_1, nx13315, 
      nx13608, nx13612, label_7_input_2, label_7_input_state_machine_2, 
      nx13640, nx13644, nx13662, label_7_input_3, 
      label_7_input_state_machine_3, nx13319, nx13672, nx13676, 
      label_7_input_4, label_7_input_state_machine_4, nx13704, nx13708, 
      nx13726, label_7_input_5, label_7_input_state_machine_5, nx13321, 
      nx13736, nx13740, label_7_input_6, label_7_input_state_machine_6, 
      nx13768, nx13772, nx13790, label_7_input_7, 
      label_7_input_state_machine_7, nx13323, nx13800, nx13804, 
      label_7_input_8, label_7_input_state_machine_8, nx13832, nx13836, 
      nx13854, label_7_input_9, label_7_input_state_machine_9, nx13325, 
      nx13864, nx13868, label_7_input_10, label_7_input_state_machine_10, 
      nx13896, nx13900, nx13918, label_7_input_11, 
      label_7_input_state_machine_11, nx13329, nx13928, nx13932, 
      label_7_input_12, label_7_input_state_machine_12, nx13960, nx13964, 
      nx13982, label_7_input_13, label_7_input_state_machine_13, nx13332, 
      nx13992, nx13996, nx14018, nx14022, label_8_input_14, 
      label_8_input_state_machine_14, label_8_input_0, 
      booth_booth_integrtaion_7_shift_reg_output_9, 
      booth_booth_integrtaion_7_shift_Reg_count_9, 
      booth_booth_integrtaion_7_shift_Reg_output_8, 
      booth_booth_integrtaion_7_shift_Reg_count_8, 
      booth_booth_integrtaion_7_shift_Reg_output_7, 
      booth_booth_integrtaion_7_shift_Reg_count_7, 
      booth_booth_integrtaion_7_shift_Reg_output_6, 
      booth_booth_integrtaion_7_shift_Reg_count_6, 
      booth_booth_integrtaion_7_shift_Reg_output_5, 
      booth_booth_integrtaion_7_shift_Reg_count_5, 
      booth_booth_integrtaion_7_shift_Reg_output_4, 
      booth_booth_integrtaion_7_shift_Reg_count_4, 
      booth_booth_integrtaion_7_shift_Reg_output_3, 
      booth_booth_integrtaion_7_shift_Reg_count_3, 
      booth_booth_integrtaion_7_shift_Reg_output_2, 
      booth_booth_integrtaion_7_shift_Reg_count_2, 
      booth_booth_integrtaion_7_shift_Reg_output_1, 
      booth_booth_integrtaion_7_shift_Reg_count_1, 
      booth_booth_integrtaion_7_shift_reg_output_0, 
      booth_booth_integrtaion_7_shift_Reg_count_0, 
      booth_booth_integration_output_7_1, booth_booth_integration_output_7_2, 
      booth_booth_integration_output_7_3, booth_booth_integration_output_7_4, 
      booth_booth_integration_output_7_5, booth_booth_integration_output_7_6, 
      booth_booth_integration_output_7_7, booth_booth_integration_output_7_8, 
      booth_booth_integration_output_7_9, 
      booth_booth_integration_output_7_10, 
      booth_booth_integration_output_7_11, 
      booth_booth_integration_output_7_12, 
      booth_booth_integration_output_7_13, 
      booth_booth_integration_output_7_14, 
      booth_booth_integration_output_7_15, 
      booth_booth_integrtaion_7_booth_output_16, nx14152, nx14158, 
      booth_booth_integrtaion_7_booth_output_17, nx13334, nx14166, nx14182, 
      booth_booth_integrtaion_7_booth_output_18, nx13335, nx14192, nx14196, 
      nx14210, booth_booth_integrtaion_7_booth_output_19, nx13336, nx14216, 
      nx14220, nx14230, booth_booth_integrtaion_7_booth_output_20, nx13337, 
      nx14240, nx14244, nx14258, booth_booth_integrtaion_7_booth_output_21, 
      nx13339, nx14264, nx14268, nx14278, 
      booth_booth_integrtaion_7_booth_output_22, nx13341, nx14288, nx14292, 
      nx14306, booth_booth_integrtaion_7_booth_output_23, nx13343, nx14312, 
      nx14316, nx14326, booth_booth_integrtaion_7_booth_output_24, nx13344, 
      nx14336, nx14340, nx14354, booth_booth_integrtaion_7_booth_output_25, 
      nx13345, nx14360, nx14364, nx14374, 
      booth_booth_integrtaion_7_booth_output_26, nx13346, nx14384, nx14388, 
      nx14402, booth_booth_integrtaion_7_booth_output_27, nx13347, nx14408, 
      nx14412, nx14422, booth_booth_integrtaion_7_booth_output_28, nx13348, 
      nx14432, nx14436, nx14450, booth_booth_integrtaion_7_booth_output_29, 
      nx13349, nx14456, nx14460, nx14470, 
      booth_booth_integrtaion_7_booth_output_31, nx13351, nx14480, nx14484, 
      nx14498, nx14500, nx14508, nx14514, nx14522, nx14538, nx14546, nx14562, 
      nx14570, nx14586, nx14594, nx14610, nx14618, nx14634, nx14642, nx14658, 
      nx14666, nx14682, nx14688, nx14694, nx14712, nx14724, nx14736, nx14748, 
      nx14760, nx14772, nx14784, nx14796, nx14808, nx14820, nx14832, nx14844, 
      nx14856, nx14868, nx14880, nx14890, label_8_input_state_machine_0, 
      nx14902, label_8_input_1, label_8_input_state_machine_1, nx13355, 
      nx14924, nx14928, label_8_input_2, label_8_input_state_machine_2, 
      nx14956, nx14960, nx14978, label_8_input_3, 
      label_8_input_state_machine_3, nx13357, nx14988, nx14992, 
      label_8_input_4, label_8_input_state_machine_4, nx15020, nx15024, 
      nx15042, label_8_input_5, label_8_input_state_machine_5, nx13359, 
      nx15052, nx15056, label_8_input_6, label_8_input_state_machine_6, 
      nx15084, nx15088, nx15106, label_8_input_7, 
      label_8_input_state_machine_7, nx13361, nx15116, nx15120, 
      label_8_input_8, label_8_input_state_machine_8, nx15148, nx15152, 
      nx15170, label_8_input_9, label_8_input_state_machine_9, nx13365, 
      nx15180, nx15184, label_8_input_10, label_8_input_state_machine_10, 
      nx15212, nx15216, nx15234, label_8_input_11, 
      label_8_input_state_machine_11, nx13368, nx15244, nx15248, 
      label_8_input_12, label_8_input_state_machine_12, nx15276, nx15280, 
      nx15298, label_8_input_13, label_8_input_state_machine_13, nx13370, 
      nx15308, nx15312, nx15334, nx15338, nx15360, 
      max_calc_comparator_fourth_inp2_13, max_calc_comparator_fourth_inp1_13, 
      max_calc_comparator_fourth_inp1_12, nx15404, 
      max_calc_comparator_fourth_inp2_11, max_calc_comparator_fourth_inp1_11, 
      max_calc_comparator_fourth_inp1_10, nx15448, 
      max_calc_comparator_fourth_inp2_9, max_calc_comparator_fourth_inp1_9, 
      max_calc_comparator_fourth_inp1_8, nx15492, 
      max_calc_comparator_fourth_inp2_7, max_calc_comparator_fourth_inp1_7, 
      max_calc_comparator_fourth_inp1_6, nx15536, 
      max_calc_comparator_fourth_inp2_5, max_calc_comparator_fourth_inp1_5, 
      max_calc_comparator_fourth_inp1_4, nx15580, 
      max_calc_comparator_fourth_inp2_3, max_calc_comparator_fourth_inp1_3, 
      max_calc_comparator_fourth_inp1_2, nx15624, 
      max_calc_comparator_fourth_inp2_1, nx15646, 
      max_calc_comparator_fourth_inp1_0, nx15682, nx15698, nx15714, nx15730, 
      nx15746, nx15762, nx15778, label_8_input_15, 
      label_8_input_state_machine_15, nx15800, nx15804, nx15808, 
      label_7_input_15, label_7_input_state_machine_15, nx15842, nx15846, 
      nx15850, nx15872, nx15874, nx15896, nx15908, 
      max_calc_comparator_second_inp2_13, max_calc_ans4_13, nx15934, 
      max_calc_comparator_second_inp1_13, max_calc_ans3_13, nx15970, 
      max_calc_ans4_12, nx16008, max_calc_comparator_second_inp1_12, 
      max_calc_ans3_12, nx16044, nx16056, max_calc_comparator_second_inp2_11, 
      max_calc_ans4_11, nx16082, max_calc_comparator_second_inp1_11, 
      max_calc_ans3_11, nx16118, max_calc_ans4_10, nx16156, 
      max_calc_comparator_second_inp1_10, max_calc_ans3_10, nx16192, nx16204, 
      max_calc_comparator_second_inp2_9, max_calc_ans4_9, nx16230, 
      max_calc_comparator_second_inp1_9, max_calc_ans3_9, nx16266, 
      max_calc_ans4_8, nx16304, max_calc_comparator_second_inp1_8, 
      max_calc_ans3_8, nx16340, nx16352, max_calc_comparator_second_inp2_7, 
      max_calc_ans4_7, nx16378, max_calc_comparator_second_inp1_7, 
      max_calc_ans3_7, nx16414, max_calc_ans4_6, nx16452, 
      max_calc_comparator_second_inp1_6, max_calc_ans3_6, nx16488, nx16500, 
      max_calc_comparator_second_inp2_5, max_calc_ans4_5, nx16526, 
      max_calc_comparator_second_inp1_5, max_calc_ans3_5, nx16562, 
      max_calc_ans4_4, nx16600, max_calc_comparator_second_inp1_4, 
      max_calc_ans3_4, nx16636, nx16648, max_calc_comparator_second_inp2_3, 
      max_calc_ans4_3, nx16674, max_calc_comparator_second_inp1_3, 
      max_calc_ans3_3, nx16710, max_calc_ans4_2, nx16748, 
      max_calc_comparator_second_inp1_2, max_calc_ans3_2, nx16784, nx16796, 
      max_calc_comparator_second_inp2_1, max_calc_ans4_1, nx16822, 
      max_calc_ans3_1, nx16858, nx16870, max_calc_ans4_0, nx16896, 
      max_calc_comparator_second_inp1_0, max_calc_ans3_0, nx16932, nx16958, 
      nx16974, nx16990, nx17006, nx17022, nx17038, nx17054, max_calc_ans4_15, 
      nx17088, max_calc_ans3_15, nx17124, nx17136, nx17138, nx17146, nx17156, 
      max_calc_ans8_14, max_calc_comparator_first_inp1_14, max_calc_ans1_14, 
      nx13371, nx17174, max_calc_ans6_14, max_calc_ans5_14, nx17196, nx17206, 
      nx17210, nx13373, max_calc_ans7_14, nx17244, nx17248, nx17256, 
      max_calc_comparator_first_inp2_13, max_calc_ans2_13, nx17268, nx17278, 
      max_calc_ans8_13, max_calc_comparator_first_inp1_13, max_calc_ans1_13, 
      nx13375, nx17296, max_calc_ans6_13, max_calc_ans5_13, nx17318, nx17328, 
      nx17332, max_calc_ans7_13, nx17366, nx17370, 
      max_calc_comparator_first_inp2_12, max_calc_ans2_12, nx17390, nx17400, 
      max_calc_ans8_12, max_calc_comparator_first_inp1_12, max_calc_ans1_12, 
      nx13376, nx17418, max_calc_ans6_12, max_calc_ans5_12, nx17440, nx17450, 
      nx17454, max_calc_ans7_12, nx17488, nx17492, nx17500, 
      max_calc_comparator_first_inp2_11, max_calc_ans2_11, nx17512, nx17522, 
      max_calc_ans8_11, max_calc_comparator_first_inp1_11, max_calc_ans1_11, 
      nx13377, nx17540, max_calc_ans6_11, max_calc_ans5_11, nx17562, nx17572, 
      nx17576, max_calc_ans7_11, nx17610, nx17614, 
      max_calc_comparator_first_inp2_10, max_calc_ans2_10, nx17634, nx17644, 
      max_calc_ans8_10, max_calc_comparator_first_inp1_10, max_calc_ans1_10, 
      nx13379, nx17662, max_calc_ans6_10, max_calc_ans5_10, nx17684, nx17694, 
      nx17698, max_calc_ans7_10, nx17732, nx17736, nx17744, 
      max_calc_comparator_first_inp2_9, max_calc_ans2_9, nx17756, nx17766, 
      max_calc_ans8_9, max_calc_comparator_first_inp1_9, max_calc_ans1_9, 
      nx13381, nx17784, max_calc_ans6_9, max_calc_ans5_9, nx17806, nx17816, 
      nx17820, max_calc_ans7_9, nx17854, nx17858, 
      max_calc_comparator_first_inp2_8, max_calc_ans2_8, nx17878, nx17888, 
      max_calc_ans8_8, max_calc_comparator_first_inp1_8, max_calc_ans1_8, 
      nx13383, nx17906, max_calc_ans6_8, max_calc_ans5_8, nx17928, nx17938, 
      nx17942, max_calc_ans7_8, nx17976, nx17980, nx17988, 
      max_calc_comparator_first_inp2_7, max_calc_ans2_7, nx18000, nx18010, 
      max_calc_ans8_7, max_calc_comparator_first_inp1_7, max_calc_ans1_7, 
      nx13385, nx18028, max_calc_ans6_7, max_calc_ans5_7, nx18050, nx18060, 
      nx18064, max_calc_ans7_7, nx18098, nx18102, 
      max_calc_comparator_first_inp2_6, max_calc_ans2_6, nx18122, nx18132, 
      max_calc_ans8_6, max_calc_comparator_first_inp1_6, max_calc_ans1_6, 
      nx13386, nx18150, max_calc_ans6_6, max_calc_ans5_6, nx18172, nx18182, 
      nx18186, max_calc_ans7_6, nx18220, nx18224, nx18232, 
      max_calc_comparator_first_inp2_5, max_calc_ans2_5, nx18244, nx18254, 
      max_calc_ans8_5, max_calc_comparator_first_inp1_5, max_calc_ans1_5, 
      nx13387, nx18272, max_calc_ans6_5, max_calc_ans5_5, nx18294, nx18304, 
      nx18308, max_calc_ans7_5, nx18342, nx18346, 
      max_calc_comparator_first_inp2_4, max_calc_ans2_4, nx18366, nx18376, 
      max_calc_ans8_4, max_calc_comparator_first_inp1_4, max_calc_ans1_4, 
      nx13388, nx18394, max_calc_ans6_4, max_calc_ans5_4, nx18416, nx18426, 
      nx18430, max_calc_ans7_4, nx18464, nx18468, nx18476, 
      max_calc_comparator_first_inp2_3, max_calc_ans2_3, nx18488, nx18498, 
      max_calc_ans8_3, max_calc_comparator_first_inp1_3, max_calc_ans1_3, 
      nx13389, nx18516, max_calc_ans6_3, max_calc_ans5_3, nx18538, nx18548, 
      nx18552, max_calc_ans7_3, nx18586, nx18590, 
      max_calc_comparator_first_inp2_2, max_calc_ans2_2, nx18610, nx18620, 
      max_calc_ans8_2, max_calc_comparator_first_inp1_2, max_calc_ans1_2, 
      nx13391, nx18638, max_calc_ans6_2, max_calc_ans5_2, nx18660, nx18670, 
      nx18674, max_calc_ans7_2, nx18708, nx18712, nx18720, 
      max_calc_comparator_first_inp2_1, max_calc_ans2_1, nx18732, nx18742, 
      max_calc_ans8_1, max_calc_comparator_first_inp1_1, max_calc_ans1_1, 
      nx13393, nx18760, max_calc_ans6_1, max_calc_ans5_1, nx18782, nx18792, 
      nx18796, max_calc_ans7_1, nx18830, nx18834, nx18842, 
      max_calc_comparator_first_inp2_0, max_calc_ans2_0, nx18854, nx18864, 
      max_calc_ans8_0, max_calc_ans7_0, nx18888, nx18892, nx18914, nx18930, 
      nx18946, nx18962, nx18978, nx18994, nx19010, 
      max_calc_comparator_first_inp2_15, max_calc_ans2_15, nx19030, nx19040, 
      max_calc_ans8_15, max_calc_comparator_first_inp1_15, max_calc_ans1_15, 
      nx13395, nx19058, max_calc_ans6_15, max_calc_ans5_15, nx19080, nx19090, 
      nx19094, max_calc_ans7_15, nx19128, nx19132, nx19140, nx19232, nx19236, 
      nx19240, nx19250, nx19266, nx19276, nx19296, nx13403, nx13413, nx13423, 
      nx13429, nx13443, nx13453, nx13463, nx13473, nx13483, nx13493, nx13503, 
      nx13513, nx13523, nx13533, nx13543, nx13553, nx13563, nx13573, nx13583, 
      nx13593, nx13603, nx13613, nx13623, nx13633, nx13643, nx13653, nx13663, 
      nx13673, nx13683, nx13693, nx13703, nx13713, nx13723, nx13733, nx13743, 
      nx13753, nx13763, nx13773, nx13783, nx13793, nx13803, nx13813, nx13823, 
      nx13833, nx13843, nx13853, nx13863, nx13873, nx13883, nx13893, nx13903, 
      nx13913, nx13923, nx13933, nx13943, nx13953, nx13963, nx13973, nx13983, 
      nx13993, nx14003, nx14013, nx14023, nx14033, nx14043, nx14053, nx14063, 
      nx14073, nx14083, nx14093, nx14103, nx14113, nx14123, nx14133, nx14139, 
      nx14153, nx14163, nx14173, nx14183, nx14193, nx14203, nx14213, nx14223, 
      nx14233, nx14243, nx14253, nx14263, nx14273, nx14283, nx14293, nx14303, 
      nx14313, nx14323, nx14333, nx14343, nx14353, nx14363, nx14373, nx14383, 
      nx14393, nx14403, nx14413, nx14423, nx14433, nx14443, nx14453, nx14463, 
      nx14473, nx14483, nx14493, nx14503, nx14513, nx14523, nx14533, nx14543, 
      nx14553, nx14563, nx14573, nx14583, nx14593, nx14603, nx14613, nx14623, 
      nx14633, nx14643, nx14653, nx14663, nx14673, nx14683, nx14693, nx14703, 
      nx14713, nx14723, nx14733, nx14743, nx14753, nx14763, nx14773, nx14783, 
      nx14793, nx14803, nx14813, nx14823, nx14833, nx14843, nx14853, nx14863, 
      nx14873, nx14883, nx14893, nx14903, nx14913, nx14923, nx14933, nx14943, 
      nx14953, nx14963, nx14973, nx14983, nx14989, nx15003, nx15013, nx15023, 
      nx15033, nx15043, nx15053, nx15063, nx15073, nx15083, nx15093, nx15103, 
      nx15113, nx15123, nx15133, nx15143, nx15153, nx15163, nx15173, nx15183, 
      nx15193, nx15203, nx15213, nx15223, nx15233, nx15243, nx15253, nx15263, 
      nx15273, nx15283, nx15293, nx15303, nx15313, nx15323, nx15333, nx15343, 
      nx15353, nx15363, nx15373, nx15383, nx15393, nx15403, nx15413, nx15423, 
      nx15433, nx15443, nx15453, nx15463, nx15473, nx15483, nx15493, nx15503, 
      nx15513, nx15523, nx15533, nx15543, nx15553, nx15563, nx15573, nx15583, 
      nx15593, nx15603, nx15613, nx15623, nx15633, nx15643, nx15653, nx15663, 
      nx15673, nx15683, nx15693, nx15703, nx15713, nx15723, nx15733, nx15743, 
      nx15753, nx15763, nx15773, nx15783, nx15793, nx15803, nx15813, nx15823, 
      nx15833, nx15839, nx15853, nx15863, nx15873, nx15883, nx15893, nx15903, 
      nx15913, nx15923, nx15933, nx15943, nx15953, nx15963, nx15973, nx15983, 
      nx15993, nx16003, nx16013, nx16023, nx16033, nx16043, nx16053, nx16063, 
      nx16073, nx16083, nx16093, nx16103, nx16113, nx16123, nx16133, nx16143, 
      nx16153, nx16163, nx16173, nx16183, nx16193, nx16203, nx16213, nx16223, 
      nx16233, nx16243, nx16253, nx16263, nx16273, nx16283, nx16293, nx16303, 
      nx16313, nx16323, nx16333, nx16343, nx16353, nx16363, nx16373, nx16383, 
      nx16393, nx16403, nx16413, nx16423, nx16433, nx16443, nx16453, nx16463, 
      nx16473, nx16483, nx16493, nx16503, nx16513, nx16523, nx16533, nx16543, 
      nx16553, nx16563, nx16573, nx16583, nx16593, nx16603, nx16613, nx16623, 
      nx16633, nx16643, nx16653, nx16663, nx16673, nx16683, nx16689, nx16703, 
      nx16713, nx16723, nx16733, nx16743, nx16753, nx16763, nx16773, nx16783, 
      nx16793, nx16803, nx16813, nx16823, nx16833, nx16843, nx16853, nx16863, 
      nx16873, nx16883, nx16893, nx16903, nx16913, nx16923, nx16933, nx16943, 
      nx16953, nx16963, nx16973, nx16983, nx16993, nx17003, nx17013, nx17023, 
      nx17033, nx17043, nx17053, nx17063, nx17073, nx17083, nx17093, nx17103, 
      nx17113, nx17123, nx17133, nx17143, nx17153, nx17163, nx17173, nx17183, 
      nx17193, nx17203, nx17213, nx17223, nx17233, nx17243, nx17253, nx17263, 
      nx17273, nx17283, nx17293, nx17303, nx17313, nx17323, nx17333, nx17343, 
      nx17353, nx17363, nx17373, nx17383, nx17393, nx17403, nx17413, nx17423, 
      nx17433, nx17443, nx17453, nx17463, nx17473, nx17483, nx17493, nx17503, 
      nx17513, nx17523, nx17533, nx17543, nx17553, nx17563, nx17573, nx17583, 
      nx17593, nx17603, nx17609, nx17623, nx17633, nx17643, nx17653, nx17663, 
      nx17673, nx17683, nx17693, nx17703, nx17713, nx17723, nx17733, nx17743, 
      nx17753, nx17763, nx17773, nx17783, nx17793, nx17803, nx17813, nx17823, 
      nx17833, nx17843, nx17853, nx17863, nx17873, nx17883, nx17893, nx17903, 
      nx17913, nx17923, nx17933, nx17943, nx17953, nx17963, nx17973, nx17983, 
      nx17993, nx18003, nx18013, nx18023, nx18033, nx18043, nx18053, nx18063, 
      nx18073, nx18083, nx18093, nx18103, nx18113, nx18123, nx18133, nx18143, 
      nx18153, nx18163, nx18173, nx18179, nx18193, nx18203, nx18213, nx18223, 
      nx18233, nx18243, nx18253, nx18263, nx18273, nx18283, nx18293, nx18303, 
      nx18313, nx18323, nx18333, nx18343, nx18353, nx18363, nx18373, nx18383, 
      nx18393, nx18403, nx18413, nx18423, nx18433, nx18443, nx18453, nx18463, 
      nx18473, nx18483, nx18493, nx18503, nx18513, nx18523, nx18533, nx18543, 
      nx18553, nx18563, nx18573, nx18583, nx18593, nx18603, nx18613, nx18623, 
      nx18633, nx18643, nx18653, nx18663, nx18673, nx18683, nx18693, nx18703, 
      nx18713, nx18723, nx18733, nx18743, nx18753, nx18763, nx18773, nx18783, 
      nx18793, nx18803, nx18813, nx18823, nx18833, nx18843, nx18853, nx18863, 
      nx18873, nx18883, nx18893, nx18903, nx18913, nx18923, nx18933, nx18943, 
      nx18953, nx18963, nx18973, nx18983, nx18993, nx19003, nx19013, nx19023, 
      nx19033, nx19043, nx19053, nx19063, nx19073, nx19083, nx19093, nx19103, 
      nx19113, nx19123, nx19133, nx19143, nx19153, nx19163, nx19173, nx19183, 
      nx19193, nx19203, nx19213, nx19223, nx19233, nx19243, nx19253, nx19263, 
      nx19273, nx19283, nx19293, nx19303, nx19313, nx19323, nx19333, nx19343, 
      nx19353, nx19363, nx19373, nx19383, nx19393, nx19403, nx19413, nx19423, 
      nx19433, nx19443, nx19453, nx19463, nx19473, nx19483, nx19493, nx19503, 
      nx19513, nx19523, nx19533, nx19543, nx19553, nx19563, nx19573, nx19583, 
      nx19593, nx19603, nx19613, nx19623, nx19633, nx19643, nx19653, nx19659, 
      nx19673, nx19683, nx19693, nx19703, nx19713, nx19723, nx19733, nx19743, 
      nx19753, nx19763, nx19773, nx19783, nx19793, nx19803, nx19813, nx19823, 
      nx19833, nx19843, nx19853, nx19863, nx19873, nx19883, nx19893, nx19903, 
      nx19913, nx19923, nx19933, nx19943, nx19953, nx19963, nx19973, nx19983, 
      nx19993, nx20003, nx20013, nx20023, nx20033, nx20043, nx20053, nx20063, 
      nx20073, nx20083, nx20093, nx20103, nx20113, nx20123, nx20133, nx20143, 
      nx20153, nx20163, nx20173, nx20183, nx20193, nx20203, nx20213, nx20223, 
      nx20233, nx20243, nx20253, nx20263, nx20273, nx20283, nx20293, nx20303, 
      nx20313, nx20323, nx20333, nx20343, nx20353, nx20363, nx20373, nx20383, 
      nx20393, nx20403, nx20413, nx20423, nx20433, nx20443, nx20453, nx20463, 
      nx20473, nx20483, nx20493, nx20499, nx20513, nx20523, nx20533, nx20543, 
      nx20553, nx20563, nx20573, nx20583, nx20593, nx20603, nx20613, nx20623, 
      nx20633, nx20643, nx20653, nx20663, nx20673, nx20683, nx20693, nx20703, 
      nx20713, nx20723, nx20733, nx20743, nx20753, nx20763, nx20773, nx20783, 
      nx20793, nx20803, nx20813, nx20823, nx20833, nx20843, nx20853, nx20863, 
      nx20873, nx20883, nx20893, nx20903, nx20913, nx20923, nx20933, nx20943, 
      nx20953, nx20963, nx20973, nx20983, nx20993, nx21003, nx21013, nx21023, 
      nx21033, nx21043, nx21053, nx21063, nx21073, nx21083, nx21093, nx21103, 
      nx21113, nx21123, nx21133, nx21143, nx21153, nx21163, nx21173, nx21183, 
      nx21193, nx21203, nx21213, nx21223, nx21233, nx21243, nx21253, nx21263, 
      nx21273, nx21283, nx21293, nx21303, nx21313, nx21323, nx21333, nx21343, 
      nx21353, nx21363, nx21373, nx21383, nx21393, nx21403, nx21413, nx21423, 
      nx21433, nx21443, nx21453, nx21463, nx21473, nx21483, nx21493, nx21503, 
      nx21513, nx21523, nx21533, nx21543, nx21553, nx21563, nx21573, nx21583, 
      nx21593, nx21603, nx21613, nx21623, nx21633, nx21643, nx21653, nx21663, 
      nx21673, nx21683, nx21693, nx21699, nx21713, nx21723, nx21733, nx21743, 
      nx21753, nx21763, nx21773, nx21783, nx21793, nx21803, nx21813, nx21823, 
      nx21833, nx21843, nx21853, nx21863, nx21873, nx21883, nx21893, nx21903, 
      nx21913, nx21923, nx21933, nx21943, nx21953, nx21963, nx21973, nx21983, 
      nx21993, nx22003, nx22013, nx22023, nx22033, nx22043, nx22053, nx22063, 
      nx22073, nx22083, nx22093, nx22103, nx22113, nx22123, nx22133, nx22143, 
      nx22153, nx22163, nx22173, nx22183, nx22193, nx22203, nx22213, nx22223, 
      nx22233, nx22243, nx22253, nx22263, nx22273, nx22283, nx22293, nx22303, 
      nx22313, nx22323, nx22333, nx22343, nx22353, nx22363, nx22373, nx22383, 
      nx22393, nx22403, nx22413, nx22423, nx22433, nx22443, nx22453, nx22463, 
      nx22473, nx22483, nx22493, nx22503, nx22513, nx22523, nx22533, nx22539, 
      nx22553, nx22563, nx22573, nx22583, nx22593, nx22603, nx22613, nx22623, 
      nx22633, nx22643, nx22653, nx22663, nx22673, nx22683, nx22693, nx22703, 
      nx22713, nx22723, nx22733, nx22743, nx22753, nx22763, nx22773, nx22783, 
      nx22793, nx22803, nx22813, nx22823, nx22833, nx22843, nx22853, nx22863, 
      nx22873, nx22883, nx22893, nx22903, nx22913, nx22923, nx22933, nx22943, 
      nx22953, nx22963, nx22973, nx22983, nx22993, nx23003, nx23013, nx23023, 
      nx23033, nx23043, nx23053, nx23063, nx23073, nx23083, nx23093, nx23103, 
      nx23113, nx23123, nx23133, nx23143, nx23153, nx23163, nx23173, nx23183, 
      nx23193, nx23203, nx23213, nx23223, nx23233, nx23243, nx23253, nx23263, 
      nx23273, nx23283, nx23293, nx23303, nx23313, nx23323, nx23333, nx23343, 
      nx23353, nx23363, nx23373, nx23383, nx23393, nx23403, nx23413, nx23423, 
      nx23433, nx23443, nx23453, nx23463, nx23473, nx23483, nx23493, nx23503, 
      nx23513, nx23523, nx23533, nx23543, nx23553, nx23563, nx23573, nx23583, 
      nx23593, nx23603, nx23613, nx23623, nx23633, nx23643, nx23653, nx23663, 
      nx23673, nx23683, nx23693, nx23703, nx23713, nx23723, nx23733, nx23743, 
      nx23753, nx23763, nx23773, nx23783, nx23793, nx23803, nx23813, nx23823, 
      nx23833, nx23843, nx23853, nx23863, nx23873, nx23883, nx23893, nx23903, 
      nx23913, nx23923, nx23933, nx23943, nx23953, nx23963, nx23973, nx23983, 
      nx23993, nx24003, nx24013, nx24023, nx24033, nx24043, nx24053, nx24063, 
      nx24073, nx24083, nx24093, nx24103, nx24113, nx24123, nx24133, nx24143, 
      nx24153, nx24163, nx24173, nx24183, nx24193, nx24203, nx24213, nx24223, 
      nx24233, nx24243, nx24253, nx24263, nx24273, nx24283, nx24293, nx24303, 
      nx24313, nx24323, nx24333, nx24343, nx24353, nx24363, nx24373, nx24383, 
      nx24393, nx24403, nx24413, nx24423, nx24433, nx24443, nx24453, nx24463, 
      nx24473, nx24483, nx24493, nx24503, nx24513, nx24523, nx24533, nx24543, 
      nx24553, nx24563, nx24573, nx24583, nx24593, nx24603, nx24613, nx24623, 
      nx24633, nx24643, nx24653, nx24663, nx24673, nx24683, nx24693, nx24703, 
      nx24713, nx24723, nx24733, nx24743, nx24753, nx24763, nx24773, nx24783, 
      nx24793, nx24803, nx24813, nx24823, nx24833, nx24843, nx24853, nx24863, 
      nx24873, nx24883, nx24893, nx24903, nx24913, nx24923, nx24933, nx24943, 
      nx24953, nx24963, nx24973, nx24983, nx24993, nx25003, nx25013, nx25023, 
      nx25033, nx25043, nx25053, nx25063, nx25073, nx25083, nx25093, nx25103, 
      nx25113, nx25123, nx25133, nx25143, nx25153, nx25163, nx25173, nx25183, 
      nx25193, nx25203, nx25213, nx25223, nx25233, nx25243, nx25253, nx25263, 
      nx25273, nx25283, nx25293, nx25303, nx25313, nx25323, nx25333, nx25343, 
      nx25353, nx25363, nx25373, nx25383, nx25393, nx25403, nx25413, nx25423, 
      nx25433, nx25443, nx25453, nx25463, nx25473, nx25483, nx25493, nx25503, 
      nx25513, nx25523, nx25533, nx25543, nx25553, nx25563, nx25573, nx25583, 
      nx25593, nx25603, nx25613, nx25623, nx25633, nx25643, nx25653, nx25663, 
      nx25673, nx25683, nx25693, nx25703, nx25713, nx25723, nx25733, nx25743, 
      nx25753, nx25757, nx25813, nx25821, nx25823, nx25827, nx25830, nx25832, 
      nx25835, nx25849, nx25854, nx25857, nx25864, nx25874, nx25879, nx25891, 
      nx25893, nx25896, nx25900, nx25902, nx25907, nx25916, nx25919, nx25935, 
      nx25937, nx25940, nx25942, nx25944, nx25949, nx25951, nx25958, nx25962, 
      nx25975, nx25982, nx25986, nx25998, nx25999, nx26001, nx26014, nx26022, 
      nx26024, nx26027, nx26039, nx26044, nx26046, nx26052, nx26056, nx26069, 
      nx26078, nx26080, nx26083, nx26095, nx26099, nx26105, nx26109, nx26122, 
      nx26129, nx26144, nx26176, nx26180, nx26182, nx26184, nx26186, nx26188, 
      nx26191, nx26194, nx26201, nx26203, nx26223, nx26227, nx26276, nx26323, 
      nx26344, nx26349, nx26351, nx26353, nx26356, nx26360, nx26366, nx26368, 
      nx26371, nx26375, nx26381, nx26384, nx26386, nx26389, nx26391, nx26396, 
      nx26398, nx26401, nx26404, nx26412, nx26418, nx26421, nx26423, nx26426, 
      nx26428, nx26430, nx26435, nx26437, nx26440, nx26443, nx26453, nx26456, 
      nx26458, nx26461, nx26463, nx26465, nx26470, nx26472, nx26475, nx26478, 
      nx26488, nx26491, nx26493, nx26496, nx26498, nx26500, nx26505, nx26507, 
      nx26510, nx26513, nx26523, nx26526, nx26528, nx26531, nx26533, nx26535, 
      nx26540, nx26542, nx26545, nx26548, nx26558, nx26561, nx26563, nx26566, 
      nx26568, nx26570, nx26575, nx26577, nx26580, nx26583, nx26593, nx26596, 
      nx26598, nx26601, nx26603, nx26605, nx26608, nx26612, nx26615, nx26618, 
      nx26621, nx26624, nx26627, nx26630, nx26634, nx26636, nx26638, nx26640, 
      nx26642, nx26644, nx26646, nx26648, nx26661, nx26664, nx26666, nx26669, 
      nx26675, nx26693, nx26696, nx26702, nx26706, nx26755, nx26802, nx26823, 
      nx26828, nx26830, nx26832, nx26835, nx26839, nx26845, nx26847, nx26850, 
      nx26854, nx26860, nx26863, nx26865, nx26868, nx26870, nx26875, nx26877, 
      nx26880, nx26883, nx26891, nx26897, nx26900, nx26902, nx26905, nx26907, 
      nx26909, nx26914, nx26916, nx26919, nx26922, nx26932, nx26935, nx26937, 
      nx26940, nx26942, nx26944, nx26949, nx26951, nx26954, nx26957, nx26967, 
      nx26970, nx26972, nx26975, nx26977, nx26979, nx26984, nx26986, nx26989, 
      nx26992, nx27002, nx27005, nx27007, nx27010, nx27012, nx27014, nx27019, 
      nx27021, nx27024, nx27027, nx27037, nx27040, nx27042, nx27045, nx27047, 
      nx27049, nx27054, nx27056, nx27059, nx27062, nx27072, nx27075, nx27077, 
      nx27080, nx27082, nx27084, nx27087, nx27091, nx27094, nx27097, nx27100, 
      nx27103, nx27106, nx27109, nx27113, nx27115, nx27117, nx27119, nx27121, 
      nx27123, nx27125, nx27127, nx27133, nx27135, nx27141, nx27145, nx27194, 
      nx27241, nx27262, nx27267, nx27269, nx27271, nx27274, nx27278, nx27284, 
      nx27286, nx27289, nx27293, nx27299, nx27302, nx27304, nx27307, nx27309, 
      nx27314, nx27316, nx27319, nx27322, nx27330, nx27336, nx27339, nx27341, 
      nx27344, nx27346, nx27348, nx27353, nx27355, nx27358, nx27361, nx27371, 
      nx27374, nx27376, nx27379, nx27381, nx27383, nx27388, nx27390, nx27393, 
      nx27396, nx27406, nx27409, nx27411, nx27414, nx27416, nx27418, nx27423, 
      nx27425, nx27428, nx27431, nx27441, nx27444, nx27446, nx27449, nx27451, 
      nx27453, nx27458, nx27460, nx27463, nx27466, nx27476, nx27479, nx27481, 
      nx27484, nx27486, nx27488, nx27493, nx27495, nx27498, nx27501, nx27511, 
      nx27514, nx27516, nx27519, nx27521, nx27523, nx27526, nx27530, nx27533, 
      nx27536, nx27539, nx27542, nx27545, nx27548, nx27552, nx27554, nx27556, 
      nx27558, nx27560, nx27562, nx27564, nx27566, nx27571, nx27573, nx27576, 
      nx27586, nx27597, nx27608, nx27619, nx27630, nx27641, nx27652, nx27663, 
      nx27665, nx27668, nx27678, nx27679, nx27683, nx27693, nx27694, nx27698, 
      nx27708, nx27709, nx27713, nx27723, nx27724, nx27728, nx27738, nx27739, 
      nx27743, nx27753, nx27754, nx27758, nx27760, nx27763, nx27765, nx27775, 
      nx27786, nx27797, nx27808, nx27819, nx27830, nx27841, nx27852, nx27854, 
      nx27857, nx27867, nx27868, nx27872, nx27882, nx27883, nx27887, nx27897, 
      nx27898, nx27902, nx27912, nx27913, nx27917, nx27927, nx27928, nx27932, 
      nx27942, nx27943, nx27947, nx27949, nx27952, nx27956, nx27958, nx27960, 
      nx27963, nx27965, nx27967, nx27970, nx27974, nx27976, nx27980, nx27984, 
      nx27986, nx27988, nx27991, nx27993, nx27995, nx27998, nx28002, nx28004, 
      nx28008, nx28012, nx28014, nx28016, nx28019, nx28021, nx28023, nx28026, 
      nx28030, nx28032, nx28036, nx28040, nx28042, nx28044, nx28047, nx28049, 
      nx28051, nx28054, nx28058, nx28060, nx28064, nx28068, nx28070, nx28072, 
      nx28075, nx28077, nx28079, nx28082, nx28086, nx28088, nx28092, nx28096, 
      nx28098, nx28100, nx28103, nx28105, nx28107, nx28110, nx28114, nx28116, 
      nx28122, nx28124, nx28126, nx28129, nx28131, nx28137, nx28139, nx28150, 
      nx28155, nx28157, nx28168, nx28172, nx28183, nx28187, nx28236, nx28283, 
      nx28304, nx28309, nx28311, nx28313, nx28316, nx28320, nx28326, nx28328, 
      nx28331, nx28335, nx28341, nx28344, nx28346, nx28349, nx28351, nx28356, 
      nx28358, nx28361, nx28364, nx28372, nx28378, nx28381, nx28383, nx28386, 
      nx28388, nx28390, nx28395, nx28397, nx28400, nx28403, nx28413, nx28416, 
      nx28418, nx28421, nx28423, nx28425, nx28430, nx28432, nx28435, nx28438, 
      nx28448, nx28451, nx28453, nx28456, nx28458, nx28460, nx28465, nx28467, 
      nx28470, nx28473, nx28483, nx28486, nx28488, nx28491, nx28493, nx28495, 
      nx28500, nx28502, nx28505, nx28508, nx28518, nx28521, nx28523, nx28526, 
      nx28528, nx28530, nx28535, nx28537, nx28540, nx28543, nx28553, nx28556, 
      nx28558, nx28561, nx28563, nx28565, nx28568, nx28572, nx28575, nx28578, 
      nx28581, nx28584, nx28587, nx28590, nx28594, nx28596, nx28598, nx28600, 
      nx28602, nx28604, nx28606, nx28608, nx28617, nx28619, nx28626, nx28630, 
      nx28679, nx28726, nx28747, nx28752, nx28754, nx28756, nx28759, nx28763, 
      nx28769, nx28771, nx28774, nx28778, nx28784, nx28787, nx28789, nx28792, 
      nx28794, nx28799, nx28801, nx28804, nx28807, nx28815, nx28821, nx28824, 
      nx28826, nx28829, nx28831, nx28833, nx28838, nx28840, nx28843, nx28846, 
      nx28856, nx28859, nx28861, nx28864, nx28866, nx28868, nx28873, nx28875, 
      nx28878, nx28881, nx28891, nx28894, nx28896, nx28899, nx28901, nx28903, 
      nx28908, nx28910, nx28913, nx28916, nx28926, nx28929, nx28931, nx28934, 
      nx28936, nx28938, nx28943, nx28945, nx28948, nx28951, nx28961, nx28964, 
      nx28966, nx28969, nx28971, nx28973, nx28978, nx28980, nx28983, nx28986, 
      nx28996, nx28999, nx29001, nx29004, nx29006, nx29008, nx29011, nx29015, 
      nx29018, nx29021, nx29024, nx29027, nx29030, nx29033, nx29037, nx29039, 
      nx29041, nx29043, nx29045, nx29047, nx29049, nx29051, nx29061, nx29063, 
      nx29069, nx29073, nx29122, nx29169, nx29190, nx29195, nx29197, nx29199, 
      nx29202, nx29206, nx29212, nx29214, nx29217, nx29221, nx29227, nx29230, 
      nx29232, nx29235, nx29237, nx29242, nx29244, nx29247, nx29250, nx29258, 
      nx29264, nx29267, nx29269, nx29272, nx29274, nx29276, nx29281, nx29283, 
      nx29286, nx29289, nx29299, nx29302, nx29304, nx29307, nx29309, nx29311, 
      nx29316, nx29318, nx29321, nx29324, nx29334, nx29337, nx29339, nx29342, 
      nx29344, nx29346, nx29351, nx29353, nx29356, nx29359, nx29369, nx29372, 
      nx29374, nx29377, nx29379, nx29381, nx29386, nx29388, nx29391, nx29394, 
      nx29404, nx29407, nx29409, nx29412, nx29414, nx29416, nx29421, nx29423, 
      nx29426, nx29429, nx29439, nx29442, nx29444, nx29447, nx29449, nx29451, 
      nx29454, nx29458, nx29461, nx29464, nx29467, nx29470, nx29473, nx29476, 
      nx29480, nx29482, nx29484, nx29486, nx29488, nx29490, nx29492, nx29494, 
      nx29498, nx29502, nx29504, nx29510, nx29514, nx29563, nx29610, nx29631, 
      nx29636, nx29638, nx29640, nx29643, nx29647, nx29653, nx29655, nx29658, 
      nx29662, nx29668, nx29671, nx29673, nx29676, nx29678, nx29683, nx29685, 
      nx29688, nx29691, nx29699, nx29705, nx29708, nx29710, nx29713, nx29715, 
      nx29717, nx29722, nx29724, nx29727, nx29730, nx29740, nx29743, nx29745, 
      nx29748, nx29750, nx29752, nx29757, nx29759, nx29762, nx29765, nx29775, 
      nx29778, nx29780, nx29783, nx29785, nx29787, nx29792, nx29794, nx29797, 
      nx29800, nx29810, nx29813, nx29815, nx29818, nx29820, nx29822, nx29827, 
      nx29829, nx29832, nx29835, nx29845, nx29848, nx29850, nx29853, nx29855, 
      nx29857, nx29862, nx29864, nx29867, nx29870, nx29880, nx29883, nx29885, 
      nx29888, nx29890, nx29892, nx29895, nx29899, nx29902, nx29905, nx29908, 
      nx29911, nx29914, nx29917, nx29921, nx29923, nx29925, nx29927, nx29929, 
      nx29931, nx29933, nx29935, nx29940, nx29942, nx29945, nx29955, nx29966, 
      nx29977, nx29988, nx29999, nx30010, nx30021, nx30032, nx30034, nx30037, 
      nx30047, nx30048, nx30052, nx30062, nx30063, nx30067, nx30077, nx30078, 
      nx30082, nx30092, nx30093, nx30097, nx30107, nx30108, nx30112, nx30122, 
      nx30123, nx30127, nx30129, nx30132, nx30134, nx30144, nx30155, nx30166, 
      nx30177, nx30188, nx30199, nx30210, nx30221, nx30223, nx30226, nx30236, 
      nx30237, nx30241, nx30251, nx30252, nx30256, nx30266, nx30267, nx30271, 
      nx30281, nx30282, nx30286, nx30296, nx30297, nx30301, nx30311, nx30312, 
      nx30316, nx30318, nx30321, nx30325, nx30327, nx30329, nx30332, nx30334, 
      nx30336, nx30339, nx30343, nx30345, nx30349, nx30353, nx30355, nx30357, 
      nx30360, nx30362, nx30364, nx30367, nx30371, nx30373, nx30377, nx30381, 
      nx30383, nx30385, nx30388, nx30390, nx30392, nx30395, nx30399, nx30401, 
      nx30405, nx30409, nx30411, nx30413, nx30416, nx30418, nx30420, nx30423, 
      nx30427, nx30429, nx30433, nx30437, nx30439, nx30441, nx30444, nx30446, 
      nx30448, nx30451, nx30455, nx30457, nx30461, nx30465, nx30467, nx30469, 
      nx30472, nx30474, nx30476, nx30479, nx30483, nx30485, nx30491, nx30493, 
      nx30495, nx30498, nx30500, nx30506, nx30508, nx30519, nx30524, nx30526, 
      nx30537, nx30546, nx30548, nx30555, nx30559, nx30608, nx30655, nx30676, 
      nx30681, nx30683, nx30685, nx30688, nx30692, nx30698, nx30700, nx30703, 
      nx30707, nx30713, nx30716, nx30718, nx30721, nx30723, nx30728, nx30730, 
      nx30733, nx30736, nx30744, nx30750, nx30753, nx30755, nx30758, nx30760, 
      nx30762, nx30767, nx30769, nx30772, nx30775, nx30785, nx30788, nx30790, 
      nx30793, nx30795, nx30797, nx30802, nx30804, nx30807, nx30810, nx30820, 
      nx30823, nx30825, nx30828, nx30830, nx30832, nx30837, nx30839, nx30842, 
      nx30845, nx30855, nx30858, nx30860, nx30863, nx30865, nx30867, nx30872, 
      nx30874, nx30877, nx30880, nx30890, nx30893, nx30895, nx30898, nx30900, 
      nx30902, nx30907, nx30909, nx30912, nx30915, nx30925, nx30928, nx30930, 
      nx30933, nx30935, nx30937, nx30940, nx30944, nx30947, nx30950, nx30953, 
      nx30956, nx30959, nx30962, nx30966, nx30968, nx30970, nx30972, nx30974, 
      nx30976, nx30978, nx30980, nx30990, nx30992, nx30998, nx31002, nx31051, 
      nx31098, nx31119, nx31124, nx31126, nx31128, nx31131, nx31135, nx31141, 
      nx31143, nx31146, nx31150, nx31156, nx31159, nx31161, nx31164, nx31166, 
      nx31171, nx31173, nx31176, nx31179, nx31187, nx31193, nx31196, nx31198, 
      nx31201, nx31203, nx31205, nx31210, nx31212, nx31215, nx31218, nx31228, 
      nx31231, nx31233, nx31236, nx31238, nx31240, nx31245, nx31247, nx31250, 
      nx31253, nx31263, nx31266, nx31268, nx31271, nx31273, nx31275, nx31280, 
      nx31282, nx31285, nx31288, nx31298, nx31301, nx31303, nx31306, nx31308, 
      nx31310, nx31315, nx31317, nx31320, nx31323, nx31333, nx31336, nx31338, 
      nx31341, nx31343, nx31345, nx31350, nx31352, nx31355, nx31358, nx31368, 
      nx31371, nx31373, nx31376, nx31378, nx31380, nx31383, nx31387, nx31390, 
      nx31393, nx31396, nx31399, nx31402, nx31405, nx31409, nx31411, nx31413, 
      nx31415, nx31417, nx31419, nx31421, nx31423, nx31429, nx31431, nx31437, 
      nx31441, nx31490, nx31537, nx31558, nx31563, nx31565, nx31567, nx31570, 
      nx31574, nx31580, nx31582, nx31585, nx31589, nx31595, nx31598, nx31600, 
      nx31603, nx31605, nx31610, nx31612, nx31615, nx31618, nx31626, nx31632, 
      nx31635, nx31637, nx31640, nx31642, nx31644, nx31649, nx31651, nx31654, 
      nx31657, nx31667, nx31670, nx31672, nx31675, nx31677, nx31679, nx31684, 
      nx31686, nx31689, nx31692, nx31702, nx31705, nx31707, nx31710, nx31712, 
      nx31714, nx31719, nx31721, nx31724, nx31727, nx31737, nx31740, nx31742, 
      nx31745, nx31747, nx31749, nx31754, nx31756, nx31759, nx31762, nx31772, 
      nx31775, nx31777, nx31780, nx31782, nx31784, nx31789, nx31791, nx31794, 
      nx31797, nx31807, nx31810, nx31812, nx31815, nx31817, nx31819, nx31822, 
      nx31826, nx31829, nx31832, nx31835, nx31838, nx31841, nx31844, nx31848, 
      nx31850, nx31852, nx31854, nx31856, nx31858, nx31860, nx31862, nx31867, 
      nx31869, nx31872, nx31882, nx31893, nx31904, nx31915, nx31926, nx31937, 
      nx31948, nx31959, nx31961, nx31964, nx31974, nx31975, nx31979, nx31989, 
      nx31990, nx31994, nx32004, nx32005, nx32009, nx32019, nx32020, nx32024, 
      nx32034, nx32035, nx32039, nx32049, nx32050, nx32054, nx32056, nx32059, 
      nx32061, nx32071, nx32082, nx32093, nx32104, nx32115, nx32126, nx32137, 
      nx32148, nx32150, nx32153, nx32163, nx32164, nx32168, nx32178, nx32179, 
      nx32183, nx32193, nx32194, nx32198, nx32208, nx32209, nx32213, nx32223, 
      nx32224, nx32228, nx32238, nx32239, nx32243, nx32245, nx32248, nx32252, 
      nx32254, nx32256, nx32259, nx32261, nx32263, nx32266, nx32270, nx32272, 
      nx32276, nx32280, nx32282, nx32284, nx32287, nx32289, nx32291, nx32294, 
      nx32298, nx32300, nx32304, nx32308, nx32310, nx32312, nx32315, nx32317, 
      nx32319, nx32322, nx32326, nx32328, nx32332, nx32336, nx32338, nx32340, 
      nx32343, nx32345, nx32347, nx32350, nx32354, nx32356, nx32360, nx32364, 
      nx32366, nx32368, nx32371, nx32373, nx32375, nx32378, nx32382, nx32384, 
      nx32388, nx32392, nx32394, nx32396, nx32399, nx32401, nx32403, nx32406, 
      nx32410, nx32412, nx32418, nx32420, nx32422, nx32425, nx32427, nx32433, 
      nx32435, nx32446, nx32451, nx32453, nx32464, nx32470, nx32472, nx32475, 
      nx32486, nx32497, nx32508, nx32519, nx32530, nx32541, nx32552, nx32563, 
      nx32565, nx32568, nx32578, nx32579, nx32583, nx32593, nx32594, nx32598, 
      nx32608, nx32609, nx32613, nx32623, nx32624, nx32628, nx32638, nx32639, 
      nx32643, nx32653, nx32654, nx32658, nx32660, nx32665, nx32669, nx32671, 
      nx32682, nx32693, nx32704, nx32715, nx32726, nx32737, nx32748, nx32759, 
      nx32761, nx32764, nx32774, nx32775, nx32779, nx32789, nx32790, nx32794, 
      nx32804, nx32805, nx32809, nx32819, nx32820, nx32824, nx32834, nx32835, 
      nx32839, nx32849, nx32850, nx32854, nx32856, nx32861, nx32865, nx32869, 
      nx32871, nx32880, nx32883, nx32892, nx32894, nx32897, nx32904, nx32908, 
      nx32910, nx32917, nx32921, nx32925, nx32927, nx32936, nx32939, nx32948, 
      nx32950, nx32953, nx32960, nx32964, nx32966, nx32973, nx32977, nx32981, 
      nx32983, nx32992, nx32995, nx33004, nx33006, nx33009, nx33016, nx33020, 
      nx33022, nx33029, nx33033, nx33037, nx33039, nx33048, nx33051, nx33060, 
      nx33062, nx33065, nx33072, nx33076, nx33078, nx33085, nx33089, nx33093, 
      nx33095, nx33104, nx33107, nx33116, nx33118, nx33121, nx33128, nx33132, 
      nx33134, nx33141, nx33145, nx33149, nx33151, nx33160, nx33163, nx33172, 
      nx33174, nx33177, nx33184, nx33188, nx33190, nx33197, nx33203, nx33205, 
      nx33214, nx33217, nx33226, nx33232, nx33234, nx33246, nx33257, nx33259, 
      nx33271, nx33288, nx33290, nx33292, nx33305, nx33316, nx33327, nx33338, 
      nx33349, nx33360, nx33371, nx33382, nx33384, nx33387, nx33397, nx33398, 
      nx33402, nx33412, nx33413, nx33417, nx33427, nx33428, nx33432, nx33442, 
      nx33443, nx33447, nx33457, nx33458, nx33462, nx33472, nx33473, nx33477, 
      nx33479, nx33503, nx33514, nx33525, nx33536, nx33547, nx33558, nx33569, 
      nx33580, nx33582, nx33585, nx33595, nx33596, nx33600, nx33610, nx33611, 
      nx33615, nx33625, nx33626, nx33630, nx33640, nx33641, nx33645, nx33655, 
      nx33656, nx33660, nx33670, nx33671, nx33675, nx33677, nx33694, nx33726, 
      nx33729, nx33731, nx33767, nx33799, nx33802, nx33804, nx33840, nx33872, 
      nx33875, nx33877, nx33913, nx33945, nx33948, nx33950, nx33986, nx34018, 
      nx34021, nx34023, nx34059, nx34091, nx34094, nx34096, nx34162, nx34165, 
      nx34182, nx34209, nx34359, nx34365, nx34368, nx34377, nx34380, nx34389, 
      nx34391, nx34393, nx34395, nx34397, nx34399, nx34401, nx34403, nx34405, 
      nx34407, nx34409, nx34419, nx34429, nx34457, nx34459, nx34461, nx34463, 
      nx34465, nx34467, nx34469, nx34471, nx34473, nx34475, nx34477, nx34479, 
      nx34481, nx34483, nx34485, nx34487, nx34489, nx34491, nx34493, nx34495, 
      nx34499, nx34501, nx34503, nx34505, nx34507, nx34509, nx34511, nx34513, 
      nx34515, nx34517, nx34519, nx34521, nx34523, nx34525, nx34527, nx34529, 
      nx34531, nx34533, nx34535, nx34537, nx34539, nx34541, nx34543, nx34545, 
      nx34547, nx34549, nx34551, nx34553, nx34555, nx34557, nx34571, nx34579, 
      nx34581, nx34583, nx34585, nx34587, nx34589, nx34603, nx34611, nx34613, 
      nx34615, nx34617, nx34619, nx34621, nx34635, nx34643, nx34645, nx34647, 
      nx34649, nx34651, nx34653, nx34667, nx34675, nx34677, nx34679, nx34681, 
      nx34683, nx34705, nx34735, nx34737, nx34739, nx34741, nx34743, nx34745, 
      nx34747, nx34749, nx34751, nx34753, nx34755, nx34757, nx34759, nx34761, 
      nx34763, nx34765, nx34767, nx34769, nx34771, nx34773, nx34775, nx34777, 
      nx34779, nx34781, nx34783, nx34785, nx34787, nx34789, nx34791, nx34793, 
      nx34795, nx34797, nx34799, nx34801, nx34803, nx34805, nx34807, nx34809, 
      nx34811, nx34813, nx34815, nx34817, nx34819, nx34821, nx34833, nx34847, 
      nx34855, nx34857, nx34859, nx34861, nx34863, nx34865, nx34879, nx34887, 
      nx34889, nx34891, nx34893, nx34895, nx34905, nx34913, nx34925, nx34939, 
      nx34947, nx34949, nx34951, nx34953, nx34955, nx34957, nx34971, nx34979, 
      nx34981, nx34983, nx34985, nx34987, nx34997, nx35011, nx35019, nx35021, 
      nx35023, nx35025, nx35027, nx35029, nx35043, nx35051, nx35053, nx35055, 
      nx35057, nx35059, nx35095, nx35097, nx35099, nx35101, nx35103, nx35149, 
      nx35153, nx35155, nx35157, nx35159, nx35161, nx35163, nx35165, nx35167, 
      nx35169, nx35171, nx35173, nx35175, nx35177, nx35179, nx35181, nx35183, 
      nx35185, nx35187, nx35189, nx35191, nx35193, nx35195, nx35197, nx35199, 
      nx35201, nx35205, nx35207, nx35209, nx35211, nx35213, nx35215, nx35217, 
      nx35263, nx35265, nx35267, nx35269, nx35271, nx35289, nx35301, nx35303, 
      nx35305, nx35307, nx35309, nx35313, nx35315, nx35317, nx35319, nx35321, 
      nx35323, nx35325, nx35327, nx35329, nx35331, nx35333, nx35335, nx35339, 
      nx35341, nx35343, nx35345, nx35347, nx35349, nx35351, nx35361, nx35363, 
      nx35365, nx35367, nx35369, nx35371, nx35373, nx35375, nx35377, nx35379, 
      nx35381, nx35385, nx35387, nx35389, nx35391, nx35393, nx35395, nx35397, 
      nx35399, nx35401, nx35403, nx35405, nx35407, nx35411, nx35413, nx35415, 
      nx35417, nx35419, nx35421, nx35423, nx35425, nx35427, nx35429, nx35431, 
      nx35433, nx35437, nx35439, nx35441, nx35443, nx35445, nx35447, nx35449, 
      nx35453, nx35455, nx35457, nx35459, nx35461, nx35463, nx35465, nx35467, 
      nx35469, nx35473, nx35475, nx35477, nx35479, nx35481, nx35485, nx35487, 
      nx35489, nx35491, nx35493, nx35495, nx35497, nx35499, nx35501, nx35503, 
      nx35505, nx35507, nx35511, nx35513, nx35515, nx35517, nx35519, nx35521, 
      nx35523, nx35525, nx35527, nx35529, nx35531, nx35533, nx35537, nx35539, 
      nx35541, nx35543, nx35545, nx35547, nx35549, nx35551, nx35553, nx35555, 
      nx35557, nx35559, nx35563, nx35565, nx35567, nx35569, nx35571, nx35573, 
      nx35575, nx35589, nx35591, nx35593, nx35595, nx35597, nx35599, nx35601, 
      nx35603, nx35605, nx35607, nx35609, nx35615, nx35621, nx35623, nx35625, 
      nx35627, nx35629, nx35631, nx35633, nx35635, nx35637, nx35639, nx35641, 
      nx35643, nx35645, nx35647, nx35649, nx35651, nx35653, nx35655, nx35657, 
      nx35659, nx35661, nx35663, nx35665, nx35667, nx35669, nx35671, nx35673, 
      nx35675, nx35677, nx35679, nx35681, nx35683, nx35685, nx35687, nx35689, 
      nx35691, nx35693, nx35695, nx35697, nx35699, nx35701, nx35703, nx35705, 
      nx35707, nx35709, nx35711, nx35713, nx35715, nx35717, nx35719, nx35721, 
      nx35723, nx35725, nx35727, nx35729, nx35731, nx35733, nx35735, nx35737, 
      nx35739, nx35741, nx35743, nx35745, nx35747, nx35749, nx35751, nx35753, 
      nx35755, nx35757, nx35759, nx35761, nx35763, nx35765, nx35767, nx35769, 
      nx35771, nx35773, nx35775, nx35777, nx35779, nx35781, nx35783, nx35785, 
      nx35787, nx35789, nx35791, nx35793, nx35795, nx35797, nx35799, nx35801, 
      nx35803, nx35805, nx35807, nx35809, nx35811, nx35813, nx35815, nx35817, 
      nx35819, nx35821, nx35823, nx35825, nx35827, nx35829, nx35831, nx35833, 
      nx35835, nx35837, nx35839, nx35841, nx35843, nx35845, nx35847, nx35849, 
      nx35851, nx35853, nx35855, nx35857, nx35859, nx35861, nx35863, nx35865, 
      nx35867, nx35869, nx35871, nx35873, nx35875, nx35877, nx35879, nx35881, 
      nx35883, nx35885, nx35887, nx35889, nx35891, nx35893, nx35895, nx35897, 
      nx35899, nx35901, nx35903, nx35905, nx35907, nx35909, nx35911, nx35913, 
      nx35915, nx35917, nx35919, nx35921, nx35923, nx35925, nx35927, nx35929, 
      nx35931, nx35933, nx35935, nx35937, nx35939, nx35941, nx35943, nx35945, 
      nx35947, nx35949, nx35951, nx35953, nx35955, nx35957, nx35959, nx35961, 
      nx35963, nx35965, nx35967, nx35969, nx35971, nx35973, nx35975, nx35977, 
      nx35979, nx35981, nx35983, nx35985, nx35987, nx35989, nx35991, nx35993, 
      nx35995, nx35997, nx35999, nx36001, nx36003, nx36005, nx36007, nx36009, 
      nx36011, nx36013, nx36015, nx36017, nx36019, nx36021, nx36023, nx36025, 
      nx36027, nx36029, nx36031, nx36033, nx36035, nx36037, nx36039, nx36041, 
      nx36043, nx36045, nx36047, nx36049, nx36051, nx36053, nx36055, nx36057, 
      nx36059, nx36061, nx36063, nx36065, nx36067, nx36069, nx36071, nx36073, 
      nx36075, nx36077, nx36079, nx36081, nx36083, nx36085, nx36087, nx36089, 
      nx36091, nx36093, nx36095, nx36097, nx36099, nx36101, nx36103, nx36105, 
      nx36107, nx36109, nx36111, nx36113, nx36115, nx36117, nx36119, nx36121, 
      nx36123, nx36125, nx36127, nx36129, nx36131, nx36133, nx36135, nx36137, 
      nx36139, nx36141, nx36143, nx36145, nx36147, nx36149, nx36151, nx36153, 
      nx36155, nx36157, nx36159, nx36161, nx36163, nx36165, nx36167, nx36169, 
      nx36171, nx36173, nx36175, nx36177, nx36179, nx36181, nx36183, nx36185, 
      nx36187, nx36189, nx36191, nx36193, nx36195, nx36197, nx36199, nx36201, 
      nx36203, nx36205, nx36207, nx36209, nx36211, nx36213, nx36215, nx36217, 
      nx36219, nx36221, nx36223, nx36225, nx36227, nx36229, nx36231, nx36233, 
      nx36235, nx36237, nx36239, nx36241, nx36243, nx36245, nx36247, nx36249, 
      nx36251, nx36253, nx36255, nx36257, nx36259, nx36261, nx36263, nx36265, 
      nx36267, nx36269, nx36271, nx36273, nx36275, nx36277, nx36279, nx36281, 
      nx36283, nx36285, nx36287, nx36289, nx36291, nx36293, nx36295, nx36297, 
      nx36299, nx36301, nx36307, nx36309, nx36311, nx36313, nx36315, nx36317, 
      nx36319, nx36321, nx36323, nx36325, nx36327, nx36329, nx36331, nx36333, 
      nx36335, nx36337, nx36339, nx36341, nx36343, nx36345, nx36347, nx36349, 
      nx36351, nx36353, nx36355, nx36357, nx36359, nx36361, nx36363, nx36365, 
      nx36367, nx36369, nx36371, nx36373, nx36375, nx36377, nx36379, nx36381, 
      nx36383, nx36385, nx36387, nx36389, nx36391, nx36393: std_logic ;

begin
   enable_write <= initiate ;
   answer(15) <= answer_15_EXMPLR ;
   answer(14) <= answer_14_EXMPLR ;
   answer(13) <= answer_13_EXMPLR ;
   answer(12) <= answer_12_EXMPLR ;
   answer(11) <= answer_11_EXMPLR ;
   answer(10) <= answer_10_EXMPLR ;
   answer(9) <= answer_9_EXMPLR ;
   answer(8) <= answer_8_EXMPLR ;
   answer(7) <= answer_7_EXMPLR ;
   answer(6) <= answer_6_EXMPLR ;
   answer(5) <= answer_5_EXMPLR ;
   answer(4) <= answer_4_EXMPLR ;
   answer(3) <= answer_3_EXMPLR ;
   answer(2) <= answer_2_EXMPLR ;
   answer(1) <= answer_1_EXMPLR ;
   answer(0) <= answer_0_EXMPLR ;
   ix25758 : fake_vcc port map ( Y=>nx25757);
   booth_shift_Reg_adder_0_reg_count_18 : dffr port map ( Q=>
      enable_decoder_dst_booth, QB=>OPEN, D=>nx13613, CLK=>clk, R=>nx34461);
   booth_shift_Reg_adder_0_reg_count_17 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_17, QB=>OPEN, D=>nx13603, CLK=>clk, R=>
      nx34461);
   booth_shift_Reg_adder_0_reg_count_16 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_16, QB=>OPEN, D=>nx13593, CLK=>clk, R=>
      nx34461);
   booth_shift_Reg_adder_0_reg_count_15 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_15, QB=>OPEN, D=>nx13583, CLK=>clk, R=>
      nx34461);
   booth_shift_Reg_adder_0_reg_count_14 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_14, QB=>OPEN, D=>nx13573, CLK=>clk, R=>
      nx34461);
   booth_shift_Reg_adder_0_reg_count_13 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_13, QB=>OPEN, D=>nx13563, CLK=>clk, R=>
      nx34461);
   booth_shift_Reg_adder_0_reg_count_12 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_12, QB=>OPEN, D=>nx13553, CLK=>clk, R=>
      nx34459);
   booth_shift_Reg_adder_0_reg_count_11 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_11, QB=>OPEN, D=>nx13543, CLK=>clk, R=>
      nx34459);
   booth_shift_Reg_adder_0_reg_count_10 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_10, QB=>OPEN, D=>nx13533, CLK=>clk, R=>
      nx34459);
   booth_shift_Reg_adder_0_reg_count_9 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_9, QB=>OPEN, D=>nx13523, CLK=>clk, R=>
      nx34459);
   booth_shift_Reg_adder_0_reg_count_8 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_8, QB=>OPEN, D=>nx13513, CLK=>clk, R=>
      nx34459);
   booth_shift_Reg_adder_0_reg_count_7 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_7, QB=>OPEN, D=>nx13503, CLK=>clk, R=>
      nx34459);
   booth_shift_Reg_adder_0_reg_count_6 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_6, QB=>OPEN, D=>nx13493, CLK=>clk, R=>
      nx34459);
   booth_shift_Reg_adder_0_reg_count_5 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_5, QB=>OPEN, D=>nx13483, CLK=>clk, R=>
      nx35615);
   booth_shift_Reg_adder_0_reg_count_4 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_4, QB=>OPEN, D=>nx13473, CLK=>clk, R=>
      nx35615);
   booth_shift_Reg_adder_0_reg_count_3 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_3, QB=>OPEN, D=>nx13463, CLK=>clk, R=>
      nx35615);
   booth_shift_Reg_adder_0_reg_count_2 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_2, QB=>OPEN, D=>nx13453, CLK=>clk, R=>
      nx35615);
   booth_shift_Reg_adder_0_reg_count_1 : dffr port map ( Q=>
      booth_shift_Reg_adder_0_output_1, QB=>OPEN, D=>nx13443, CLK=>clk, R=>
      nx35615);
   booth_shift_Reg_adder_0_reg_count_0 : dffs_ni port map ( Q=>
      booth_shift_Reg_adder_0_output_0, QB=>OPEN, D=>nx13429, CLK=>clk, S=>
      nx35615);
   reg_ready_signal : dffr port map ( Q=>ready_signal, QB=>OPEN, D=>nx13423, 
      CLK=>clk, R=>rst);
   ix14104 : mux21_ni port map ( Y=>nx14103, A0=>state(0), A1=>nx830, S0=>
      nx12877);
   ix517 : nor03_2x port map ( Y=>nx516, A0=>num_out_2, A1=>num_out_0, A2=>
      num_out_1);
   num_loop1_2_fx_reg_q : dffr port map ( Q=>num_out_2, QB=>OPEN, D=>nx13833, 
      CLK=>clk, R=>rst);
   reg_num_in_2 : dff port map ( Q=>num_in_2, QB=>OPEN, D=>nx13823, CLK=>clk
   );
   ix13824 : mux21_ni port map ( Y=>nx13823, A0=>nx496, A1=>num_in_2, S0=>
      nx35161);
   ix25822 : xnor2 port map ( Y=>nx25821, A0=>nx25823, A1=>nx25986);
   ix25824 : aoi22 port map ( Y=>nx25823, A0=>nx34501, A1=>alu_inp1_1, B0=>
      nx412, B1=>nx12898);
   ix25828 : nand03 port map ( Y=>nx25827, A0=>nx278, A1=>nx25940, A2=>
      nx26129);
   ix279 : nand02 port map ( Y=>nx278, A0=>nx25830, A1=>nx12887);
   ix25831 : aoi32 port map ( Y=>nx25830, A0=>nx25832, A1=>nx12882, A2=>
      nx266, B0=>nx25900, B1=>nx258);
   ix25833 : nand02 port map ( Y=>nx25832, A0=>nx12891, A1=>nx12879);
   ix789 : nor04_2x port map ( Y=>nx12891, A0=>nx25835, A1=>num_out_3, A2=>
      num_out_4, A3=>nx26044);
   num_loop1_0_fx_reg_q : dffr port map ( Q=>num_out_0, QB=>OPEN, D=>nx13713, 
      CLK=>clk, R=>rst);
   reg_num_in_0 : dff port map ( Q=>num_in_0, QB=>OPEN, D=>nx13703, CLK=>clk
   );
   ix13704 : mux21_ni port map ( Y=>nx13703, A0=>nx376, A1=>num_in_0, S0=>
      nx35159);
   ix13644 : mux21_ni port map ( Y=>nx13643, A0=>nx34393, A1=>nx210, S0=>
      nx12877);
   ix211 : nand03 port map ( Y=>nx210, A0=>nx25849, A1=>nx35103, A2=>nx35149
   );
   ix25850 : nand02 port map ( Y=>nx25849, A0=>nx25813, A1=>nx12879);
   reg_state_1 : dffr port map ( Q=>state(1), QB=>OPEN, D=>nx13643, CLK=>clk, 
      R=>rst);
   ix25855 : nand02 port map ( Y=>nx25854, A0=>nx34397, A1=>nx172);
   reg_state_0 : dffr port map ( Q=>state(0), QB=>nx25857, D=>nx14103, CLK=>
      clk, R=>rst);
   reg_state_2 : dffr port map ( Q=>state(2), QB=>OPEN, D=>nx14093, CLK=>clk, 
      R=>rst);
   reg_alu_inp1_0 : dff port map ( Q=>alu_inp1_0, QB=>OPEN, D=>nx13723, CLK
      =>clk);
   ix13724 : mux21_ni port map ( Y=>nx13723, A0=>nx390, A1=>alu_inp1_0, S0=>
      nx35095);
   address_loop1_0_fx_reg_q : dffr port map ( Q=>address_out_0, QB=>OPEN, D
      =>nx13693, CLK=>clk, R=>rst);
   ix13694 : mux21_ni port map ( Y=>nx13693, A0=>address_out_0, A1=>
      address_in_0, S0=>nx34503);
   reg_address_in_0 : dffr port map ( Q=>address_in_0, QB=>OPEN, D=>nx13683, 
      CLK=>clk, R=>rst);
   ix13684 : mux21_ni port map ( Y=>nx13683, A0=>address_in_0, A1=>nx358, S0
      =>nx34507);
   ix359 : nor02_2x port map ( Y=>nx358, A0=>nx25864, A1=>nx35787);
   reg_sub_state_1 : dffr port map ( Q=>sub_state(1), QB=>OPEN, D=>nx13413, 
      CLK=>clk, R=>rst);
   ix13414 : mux21_ni port map ( Y=>nx13413, A0=>sub_state(1), A1=>nx26, S0
      =>nx12883);
   ix25880 : oai21 port map ( Y=>nx25879, A0=>sub_state(1), A1=>nx34401, B0
      =>nx35157);
   reg_sub_state_0 : dffr port map ( Q=>sub_state(0), QB=>OPEN, D=>nx13403, 
      CLK=>clk, R=>rst);
   ix13404 : mux21_ni port map ( Y=>nx13403, A0=>nx34401, A1=>nx20, S0=>
      nx12883);
   ix183 : oai22 port map ( Y=>nx12883, A0=>nx35155, A1=>nx25891, B0=>
      nx12879, B1=>nx25893);
   ix25892 : nand02 port map ( Y=>nx25891, A0=>nx25813, A1=>nx12879);
   ix25897 : aoi21 port map ( Y=>nx25896, A0=>sub_state(1), A1=>nx34401, B0
      =>nx34397);
   ix351 : oai43 port map ( Y=>nx350, A0=>nx35155, A1=>nx12891, A2=>nx25900, 
      A3=>nx25902, B0=>nx25919, B1=>nx34389, B2=>nx34393);
   ix25903 : oai21 port map ( Y=>nx25902, A0=>nx334, A1=>nx25916, B0=>nx258
   );
   ix259 : nor02_2x port map ( Y=>nx258, A0=>nx34401, A1=>nx25879);
   reg_sub_state_2 : dffr port map ( Q=>sub_state(2), QB=>OPEN, D=>nx13633, 
      CLK=>clk, R=>rst);
   ix321 : xnor2 port map ( Y=>nx320, A0=>sub_state(1), A1=>nx34401);
   reg_enable_address : dff port map ( Q=>enable_address, QB=>OPEN, D=>
      nx13673, CLK=>clk);
   ix13674 : or02 port map ( Y=>nx13673, A0=>nx34503, A1=>nx300);
   ix301 : nor03_2x port map ( Y=>nx300, A0=>nx38, A1=>rst, A2=>nx35099);
   ix39 : nand02 port map ( Y=>nx38, A0=>nx35157, A1=>nx34401);
   ix13734 : nand02 port map ( Y=>nx13733, A0=>nx25935, A1=>nx35095);
   reg_alu_inp2_0 : dff port map ( Q=>OPEN, QB=>nx25935, D=>nx13733, CLK=>
      clk);
   ix25938 : nand03 port map ( Y=>nx25937, A0=>nx242, A1=>nx25940, A2=>
      nx25942);
   ix25941 : inv01 port map ( Y=>nx25940, A=>rst);
   ix25943 : nand02 port map ( Y=>nx25942, A0=>nx25944, A1=>nx34405);
   ix25945 : nor03_2x port map ( Y=>nx25944, A0=>sub_state(1), A1=>nx34403, 
      A2=>nx34397);
   ix13654 : nand02 port map ( Y=>nx13653, A0=>nx35795, A1=>nx25951);
   reg_enable_num : dffr port map ( Q=>OPEN, QB=>nx25949, D=>nx13653, CLK=>
      clk, R=>rst);
   ix25952 : nand02 port map ( Y=>nx25951, A0=>nx34495, A1=>nx25944);
   num_loop1_1_fx_reg_q : dffr port map ( Q=>num_out_1, QB=>OPEN, D=>nx13773, 
      CLK=>clk, R=>rst);
   ix13764 : mux21 port map ( Y=>nx13763, A0=>nx25958, A1=>nx25975, S0=>
      nx35159);
   ix25959 : aoi22 port map ( Y=>nx25958, A0=>mdr_data_out(1), A1=>nx34495, 
      B0=>nx414, B1=>nx34405);
   ix415 : xnor2 port map ( Y=>nx414, A0=>nx412, A1=>nx25962);
   reg_alu_inp1_1 : dff port map ( Q=>alu_inp1_1, QB=>OPEN, D=>nx13783, CLK
      =>clk);
   ix13784 : mux21_ni port map ( Y=>nx13783, A0=>nx448, A1=>alu_inp1_1, S0=>
      nx35095);
   address_loop1_1_fx_reg_q : dffr port map ( Q=>address_out_1, QB=>OPEN, D
      =>nx13753, CLK=>clk, R=>rst);
   ix13754 : mux21_ni port map ( Y=>nx13753, A0=>address_out_1, A1=>
      address_in_1, S0=>nx34503);
   reg_address_in_1 : dffr port map ( Q=>address_in_1, QB=>OPEN, D=>nx13743, 
      CLK=>clk, R=>rst);
   ix13744 : mux21_ni port map ( Y=>nx13743, A0=>address_in_1, A1=>nx416, S0
      =>nx34507);
   ix417 : nor02ii port map ( Y=>nx416, A0=>nx35787, A1=>nx414);
   reg_num_in_1 : dff port map ( Q=>num_in_1, QB=>nx25975, D=>nx13763, CLK=>
      clk);
   num_loop1_3_fx_reg_q : dffr port map ( Q=>num_out_3, QB=>OPEN, D=>nx13883, 
      CLK=>clk, R=>rst);
   ix13874 : mux21 port map ( Y=>nx13873, A0=>nx25982, A1=>nx26014, S0=>
      nx35159);
   ix25983 : aoi22 port map ( Y=>nx25982, A0=>mdr_data_out(3), A1=>nx34495, 
      B0=>nx12901, B1=>nx34405);
   ix551 : xnor2 port map ( Y=>nx12901, A0=>nx522, A1=>nx26001);
   ix523 : oai22 port map ( Y=>nx522, A0=>nx25823, A1=>nx25986, B0=>nx35799, 
      B1=>nx25998);
   reg_alu_inp1_2 : dff port map ( Q=>alu_inp1_2, QB=>nx25998, D=>nx13813, 
      CLK=>clk);
   ix13814 : mux21_ni port map ( Y=>nx13813, A0=>nx480, A1=>alu_inp1_2, S0=>
      nx35095);
   address_loop1_2_fx_reg_q : dffr port map ( Q=>address_out_2, QB=>OPEN, D
      =>nx13803, CLK=>clk, R=>rst);
   ix13804 : mux21_ni port map ( Y=>nx13803, A0=>address_out_2, A1=>
      address_in_2, S0=>nx34503);
   reg_address_in_2 : dffr port map ( Q=>address_in_2, QB=>OPEN, D=>nx13793, 
      CLK=>clk, R=>rst);
   ix13794 : mux21_ni port map ( Y=>nx13793, A0=>address_in_2, A1=>nx464, S0
      =>nx34507);
   ix465 : nor02_2x port map ( Y=>nx464, A0=>nx25821, A1=>nx35787);
   reg_alu_sel : dff port map ( Q=>OPEN, QB=>nx25999, D=>nx13663, CLK=>clk);
   reg_alu_inp1_3 : dff port map ( Q=>alu_inp1_3, QB=>OPEN, D=>nx13863, CLK
      =>clk);
   ix13864 : mux21_ni port map ( Y=>nx13863, A0=>nx540, A1=>alu_inp1_3, S0=>
      nx35095);
   address_loop1_3_fx_reg_q : dffr port map ( Q=>address_out_3, QB=>OPEN, D
      =>nx13853, CLK=>clk, R=>rst);
   ix13854 : mux21_ni port map ( Y=>nx13853, A0=>address_out_3, A1=>
      address_in_3, S0=>nx34503);
   reg_address_in_3 : dffr port map ( Q=>address_in_3, QB=>OPEN, D=>nx13843, 
      CLK=>clk, R=>rst);
   ix13844 : mux21_ni port map ( Y=>nx13843, A0=>address_in_3, A1=>nx524, S0
      =>nx34507);
   ix525 : nor02ii port map ( Y=>nx524, A0=>nx35787, A1=>nx12901);
   reg_num_in_3 : dff port map ( Q=>num_in_3, QB=>nx26014, D=>nx13873, CLK=>
      clk);
   num_loop1_4_fx_reg_q : dffr port map ( Q=>num_out_4, QB=>OPEN, D=>nx13933, 
      CLK=>clk, R=>rst);
   reg_num_in_4 : dff port map ( Q=>num_in_4, QB=>OPEN, D=>nx13923, CLK=>clk
   );
   ix13924 : mux21_ni port map ( Y=>nx13923, A0=>nx606, A1=>num_in_4, S0=>
      nx35159);
   ix26023 : xnor2 port map ( Y=>nx26022, A0=>nx26024, A1=>nx26027);
   ix26025 : aoi22 port map ( Y=>nx26024, A0=>nx34499, A1=>alu_inp1_3, B0=>
      nx522, B1=>nx548);
   reg_alu_inp1_4 : dff port map ( Q=>alu_inp1_4, QB=>nx26039, D=>nx13913, 
      CLK=>clk);
   ix13914 : mux21_ni port map ( Y=>nx13913, A0=>nx590, A1=>alu_inp1_4, S0=>
      nx35095);
   address_loop1_4_fx_reg_q : dffr port map ( Q=>address_out_4, QB=>OPEN, D
      =>nx13903, CLK=>clk, R=>rst);
   ix13904 : mux21_ni port map ( Y=>nx13903, A0=>address_out_4, A1=>
      address_in_4, S0=>nx34503);
   reg_address_in_4 : dffr port map ( Q=>address_in_4, QB=>OPEN, D=>nx13893, 
      CLK=>clk, R=>rst);
   ix13894 : mux21_ni port map ( Y=>nx13893, A0=>address_in_4, A1=>nx574, S0
      =>nx34507);
   ix575 : nor02_2x port map ( Y=>nx574, A0=>nx26022, A1=>nx35787);
   num_loop1_5_fx_reg_q : dffr port map ( Q=>num_out_5, QB=>nx26046, D=>
      nx13983, CLK=>clk, R=>rst);
   ix13974 : mux21 port map ( Y=>nx13973, A0=>nx26052, A1=>nx26069, S0=>
      nx35159);
   ix26053 : aoi22 port map ( Y=>nx26052, A0=>mdr_data_out(5), A1=>nx34495, 
      B0=>nx12905, B1=>nx34405);
   ix659 : xnor2 port map ( Y=>nx12905, A0=>nx630, A1=>nx26056);
   ix631 : oai22 port map ( Y=>nx630, A0=>nx26024, A1=>nx26027, B0=>nx35799, 
      B1=>nx26039);
   reg_alu_inp1_5 : dff port map ( Q=>alu_inp1_5, QB=>OPEN, D=>nx13963, CLK
      =>clk);
   ix13964 : mux21_ni port map ( Y=>nx13963, A0=>nx648, A1=>alu_inp1_5, S0=>
      nx35095);
   address_loop1_5_fx_reg_q : dffr port map ( Q=>address_out_5, QB=>OPEN, D
      =>nx13953, CLK=>clk, R=>rst);
   ix13954 : mux21_ni port map ( Y=>nx13953, A0=>address_out_5, A1=>
      address_in_5, S0=>nx34503);
   reg_address_in_5 : dffr port map ( Q=>address_in_5, QB=>OPEN, D=>nx13943, 
      CLK=>clk, R=>rst);
   ix13944 : mux21_ni port map ( Y=>nx13943, A0=>address_in_5, A1=>nx632, S0
      =>nx34507);
   ix633 : nor02ii port map ( Y=>nx632, A0=>nx35787, A1=>nx12905);
   reg_num_in_5 : dff port map ( Q=>OPEN, QB=>nx26069, D=>nx13973, CLK=>clk
   );
   num_loop1_6_fx_reg_q : dffr port map ( Q=>num_out_6, QB=>OPEN, D=>nx14033, 
      CLK=>clk, R=>rst);
   reg_num_in_6 : dff port map ( Q=>num_in_6, QB=>OPEN, D=>nx14023, CLK=>clk
   );
   ix14024 : mux21_ni port map ( Y=>nx14023, A0=>nx714, A1=>num_in_6, S0=>
      nx35159);
   ix26079 : xnor2 port map ( Y=>nx26078, A0=>nx26080, A1=>nx26083);
   ix26081 : aoi22 port map ( Y=>nx26080, A0=>nx34501, A1=>alu_inp1_5, B0=>
      nx630, B1=>nx656);
   reg_alu_inp1_6 : dff port map ( Q=>alu_inp1_6, QB=>nx26095, D=>nx14013, 
      CLK=>clk);
   ix14014 : mux21_ni port map ( Y=>nx14013, A0=>nx698, A1=>alu_inp1_6, S0=>
      nx35097);
   address_loop1_6_fx_reg_q : dffr port map ( Q=>address_out_6, QB=>OPEN, D
      =>nx14003, CLK=>clk, R=>rst);
   ix14004 : mux21_ni port map ( Y=>nx14003, A0=>address_out_6, A1=>
      address_in_6, S0=>nx34505);
   reg_address_in_6 : dffr port map ( Q=>address_in_6, QB=>OPEN, D=>nx13993, 
      CLK=>clk, R=>rst);
   ix13994 : mux21_ni port map ( Y=>nx13993, A0=>address_in_6, A1=>nx682, S0
      =>nx34507);
   ix683 : nor02_2x port map ( Y=>nx682, A0=>nx26078, A1=>nx35787);
   num_loop1_7_fx_reg_q : dffr port map ( Q=>num_out_7, QB=>nx26099, D=>
      nx14083, CLK=>clk, R=>rst);
   ix14074 : mux21 port map ( Y=>nx14073, A0=>nx26105, A1=>nx26122, S0=>
      nx35159);
   ix26106 : aoi22 port map ( Y=>nx26105, A0=>mdr_data_out(7), A1=>nx34495, 
      B0=>nx12907, B1=>nx34407);
   ix765 : xnor2 port map ( Y=>nx12907, A0=>nx736, A1=>nx26109);
   ix737 : oai22 port map ( Y=>nx736, A0=>nx26080, A1=>nx26083, B0=>nx35799, 
      B1=>nx26095);
   reg_alu_inp1_7 : dff port map ( Q=>alu_inp1_7, QB=>OPEN, D=>nx14063, CLK
      =>clk);
   ix14064 : mux21_ni port map ( Y=>nx14063, A0=>nx754, A1=>alu_inp1_7, S0=>
      nx35097);
   address_loop1_7_fx_reg_q : dffr port map ( Q=>address_out_7, QB=>OPEN, D
      =>nx14053, CLK=>clk, R=>rst);
   ix14054 : mux21_ni port map ( Y=>nx14053, A0=>address_out_7, A1=>
      address_in_7, S0=>nx34505);
   reg_address_in_7 : dffr port map ( Q=>address_in_7, QB=>OPEN, D=>nx14043, 
      CLK=>clk, R=>rst);
   ix14044 : mux21_ni port map ( Y=>nx14043, A0=>address_in_7, A1=>nx738, S0
      =>nx34509);
   ix739 : nor02ii port map ( Y=>nx738, A0=>nx35789, A1=>nx12907);
   reg_num_in_7 : dff port map ( Q=>OPEN, QB=>nx26122, D=>nx14073, CLK=>clk
   );
   booth_shift_Reg_adder_0_reg_count_19 : dffr port map ( Q=>done, QB=>OPEN, 
      D=>nx13623, CLK=>clk, R=>nx35615);
   ix267 : aoi21 port map ( Y=>nx266, A0=>nx34403, A1=>nx174, B0=>nx38);
   ix807 : aoi21 port map ( Y=>nx12887, A0=>nx34395, A1=>state(0), B0=>
      nx34391);
   ix26130 : aoi21 port map ( Y=>nx26129, A0=>nx25942, A1=>nx846, B0=>
      nx12909);
   ix57 : nand02 port map ( Y=>nx56, A0=>nx26144, A1=>nx25832);
   ix26145 : oai21 port map ( Y=>nx26144, A0=>nx12885, A1=>nx35155, B0=>
      nx12879);
   ix12510 : fake_gnd port map ( Y=>initiate);
   max_calc_reg_done_comp : dffr port map ( Q=>done_comp, QB=>OPEN, D=>
      nx25723, CLK=>clk, R=>rst);
   ix25724 : or02 port map ( Y=>nx25723, A0=>done_comp, A1=>nx35741);
   ix17574 : oai32 port map ( Y=>nx17573, A0=>nx36389, A1=>start_comp, A2=>
      max_calc_start, B0=>nx26184, B1=>nx26191);
   max_calc_reg_state_2 : dffr port map ( Q=>max_calc_state_2, QB=>OPEN, D=>
      nx17573, CLK=>clk, R=>rst);
   ix17524 : nand02 port map ( Y=>nx17523, A0=>nx26176, A1=>nx25832);
   reg_start_comp : dffr port map ( Q=>start_comp, QB=>nx26176, D=>nx17523, 
      CLK=>clk, R=>rst);
   ix17534 : nand02 port map ( Y=>nx17533, A0=>nx26180, A1=>nx26182);
   max_calc_reg_start : dffr port map ( Q=>max_calc_start, QB=>nx26180, D=>
      nx17533, CLK=>clk, R=>rst);
   ix26185 : aoi43 port map ( Y=>nx26184, A0=>nx26186, A1=>nx34705, A2=>
      nx36389, A3=>nx26203, B0=>nx34737, B1=>nx26182, B2=>nx26201);
   ix26187 : aoi21 port map ( Y=>nx26186, A0=>nx26188, A1=>nx6300, B0=>
      nx6244);
   max_calc_reg_state_0 : dffr port map ( Q=>max_calc_state_0, QB=>nx26188, 
      D=>nx17543, CLK=>clk, R=>rst);
   ix17544 : oai32 port map ( Y=>nx17543, A0=>nx26188, A1=>start_comp, A2=>
      max_calc_start, B0=>nx26186, B1=>nx26191);
   ix6301 : aoi21 port map ( Y=>nx6300, A0=>nx36389, A1=>nx26194, B0=>
      max_calc_state_3);
   max_calc_reg_state_3 : dffr port map ( Q=>max_calc_state_3, QB=>nx26203, 
      D=>nx17563, CLK=>clk, R=>rst);
   max_calc_reg_state_1 : dffr port map ( Q=>max_calc_state_1, QB=>OPEN, D=>
      nx17553, CLK=>clk, R=>rst);
   max_calc_reg_answer_0 : dffr port map ( Q=>answer_0_EXMPLR, QB=>OPEN, D=>
      nx25563, CLK=>clk, R=>rst);
   max_calc_reg_comparator_first_inp1_0 : dff port map ( Q=>
      max_calc_comparator_first_inp1_0, QB=>OPEN, D=>nx19633, CLK=>clk);
   labelsregfile_label1_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_1_output(0), QB=>OPEN, D=>nx17223, CLK=>clk, R=>rst);
   lat_label_1_input_0 : latch port map ( Q=>label_1_input_0, D=>nx5758, CLK
      =>nx34511);
   ix5759 : oai21 port map ( Y=>nx5758, A0=>nx26223, A1=>nx34409, B0=>
      nx26227);
   reg_label_1_input_state_machine_0 : dffr port map ( Q=>
      label_1_input_state_machine_0, QB=>nx26223, D=>nx17213, CLK=>clk, R=>
      rst);
   ix26228 : oai21 port map ( Y=>nx26227, A0=>nx35731, A1=>label_1_output(0), 
      B0=>nx5746);
   booth_booth_integrtaion_0_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_1, QB=>OPEN, D=>nx17193, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_2, QB=>nx26648, D=>nx17183, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_3, QB=>OPEN, D=>nx17173, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_4, QB=>nx26646, D=>nx17163, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_5, QB=>OPEN, D=>nx17153, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_6, QB=>nx26644, D=>nx17143, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_7, QB=>OPEN, D=>nx17133, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_8, QB=>nx26642, D=>nx17123, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_9, QB=>OPEN, D=>nx17113, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_10, QB=>nx26640, D=>nx17103, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_11, QB=>OPEN, D=>nx17093, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_12, QB=>nx26638, D=>nx17083, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_13, QB=>OPEN, D=>nx17073, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_14, QB=>nx26636, D=>nx17063, CLK=>clk, 
      R=>rst);
   ix26277 : aoi22 port map ( Y=>nx26276, A0=>mdr_data_out(15), A1=>nx34667, 
      B0=>nx5544, B1=>nx5550);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_reg_output_0, QB=>OPEN, 
      D=>nx16703, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_0, QB=>OPEN, D=>nx16689, CLK
      =>clk, S=>nx34465);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_reg_output_9, QB=>OPEN, 
      D=>nx16883, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_9, QB=>OPEN, D=>nx16873, CLK
      =>clk, R=>nx34465);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_8, QB=>OPEN, 
      D=>nx16863, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_8, QB=>OPEN, D=>nx16853, CLK
      =>clk, R=>nx34465);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_7, QB=>OPEN, 
      D=>nx16843, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_7, QB=>OPEN, D=>nx16833, CLK
      =>clk, R=>nx34463);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_6, QB=>OPEN, 
      D=>nx16823, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_6, QB=>OPEN, D=>nx16813, CLK
      =>clk, R=>nx34463);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_5, QB=>OPEN, 
      D=>nx16803, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_5, QB=>OPEN, D=>nx16793, CLK
      =>clk, R=>nx34463);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_4, QB=>OPEN, 
      D=>nx16783, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_4, QB=>OPEN, D=>nx16773, CLK
      =>clk, R=>nx34463);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_3, QB=>OPEN, 
      D=>nx16763, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_3, QB=>OPEN, D=>nx16753, CLK
      =>clk, R=>nx34463);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_2, QB=>OPEN, 
      D=>nx16743, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_2, QB=>OPEN, D=>nx16733, CLK
      =>clk, R=>nx34463);
   booth_booth_integrtaion_0_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_0_shift_Reg_output_1, QB=>OPEN, 
      D=>nx16723, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_0_shift_Reg_count_1, QB=>OPEN, D=>nx16713, CLK
      =>clk, R=>nx34461);
   ix16684 : nand02 port map ( Y=>nx16683, A0=>nx35803, A1=>nx34653);
   booth_booth_integrtaion_0_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx26323, D=>nx16683, CLK=>clk, S=>nx34463);
   ix5545 : nand02 port map ( Y=>nx5544, A0=>nx26344, A1=>nx26356);
   ix26345 : oai21 port map ( Y=>nx26344, A0=>nx34681, A1=>nx34675, B0=>
      mdr_data_out(16));
   ix16894 : oai21 port map ( Y=>nx16893, A0=>nx26349, A1=>nx35193, B0=>
      nx26351);
   booth_booth_integrtaion_0_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx26349, D=>nx16893, CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx26353, D=>nx17203, CLK=>clk, R=>rst);
   ix26361 : xnor2 port map ( Y=>nx26360, A0=>nx5014, A1=>nx13067);
   ix17034 : oai21 port map ( Y=>nx17033, A0=>nx26366, A1=>nx35193, B0=>
      nx26368);
   booth_booth_integrtaion_0_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_17, QB=>nx26366, D=>nx17033, 
      CLK=>clk, R=>rst);
   ix26369 : nand03 port map ( Y=>nx26368, A0=>nx35201, A1=>nx5522, A2=>
      nx36003);
   ix5523 : xnor2 port map ( Y=>nx5522, A0=>nx26371, A1=>nx13069);
   ix26372 : aoi22 port map ( Y=>nx26371, A0=>
      booth_booth_integrtaion_0_booth_output_17, A1=>nx5038, B0=>nx5014, B1
      =>nx13067);
   ix5023 : nand02 port map ( Y=>nx5022, A0=>mdr_data_out(17), A1=>
      mdr_data_out(16));
   ix26376 : or02 port map ( Y=>nx26375, A0=>mdr_data_out(16), A1=>
      mdr_data_out(17));
   ix26382 : xnor2 port map ( Y=>nx26381, A0=>nx5066, A1=>nx13071);
   ix5067 : oai22 port map ( Y=>nx5066, A0=>nx26371, A1=>nx26384, B0=>
      nx26391, B1=>nx35205);
   ix26387 : aoi32 port map ( Y=>nx26386, A0=>nx5048, A1=>nx34681, A2=>
      nx26389, B0=>mdr_data_out(18), B1=>nx34675);
   ix5049 : oai21 port map ( Y=>nx5048, A0=>mdr_data_out(16), A1=>
      mdr_data_out(17), B0=>mdr_data_out(18));
   booth_booth_integrtaion_0_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_18, QB=>nx26391, D=>nx17023, 
      CLK=>clk, R=>rst);
   ix17014 : oai21 port map ( Y=>nx17013, A0=>nx26396, A1=>nx35193, B0=>
      nx26398);
   booth_booth_integrtaion_0_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_19, QB=>nx26396, D=>nx17013, 
      CLK=>clk, R=>rst);
   ix26399 : nand03 port map ( Y=>nx26398, A0=>nx35201, A1=>nx5498, A2=>
      nx36003);
   ix5499 : xnor2 port map ( Y=>nx5498, A0=>nx26401, A1=>nx13073);
   ix26402 : aoi22 port map ( Y=>nx26401, A0=>
      booth_booth_integrtaion_0_booth_output_19, A1=>nx5086, B0=>nx5066, B1
      =>nx13071);
   ix26405 : nor02ii port map ( Y=>nx26404, A0=>nx5052, A1=>mdr_data_out(19)
   );
   ix5053 : nor03_2x port map ( Y=>nx5052, A0=>mdr_data_out(18), A1=>
      mdr_data_out(16), A2=>mdr_data_out(17));
   ix5077 : nor04 port map ( Y=>nx5076, A0=>mdr_data_out(19), A1=>
      mdr_data_out(18), A2=>mdr_data_out(16), A3=>mdr_data_out(17));
   ix26419 : xnor2 port map ( Y=>nx26418, A0=>nx5114, A1=>nx13074);
   ix5115 : oai22 port map ( Y=>nx5114, A0=>nx26401, A1=>nx26421, B0=>
      nx26430, B1=>nx35207);
   ix26424 : aoi32 port map ( Y=>nx26423, A0=>nx5096, A1=>nx34681, A2=>
      nx26428, B0=>mdr_data_out(20), B1=>nx34675);
   ix5097 : nand02 port map ( Y=>nx5096, A0=>nx26426, A1=>mdr_data_out(20));
   booth_booth_integrtaion_0_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_20, QB=>nx26430, D=>nx17003, 
      CLK=>clk, R=>rst);
   ix16994 : oai21 port map ( Y=>nx16993, A0=>nx26435, A1=>nx35193, B0=>
      nx26437);
   booth_booth_integrtaion_0_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_21, QB=>nx26435, D=>nx16993, 
      CLK=>clk, R=>rst);
   ix26438 : nand03 port map ( Y=>nx26437, A0=>nx35201, A1=>nx5474, A2=>
      nx36003);
   ix5475 : xnor2 port map ( Y=>nx5474, A0=>nx26440, A1=>nx13075);
   ix26441 : aoi22 port map ( Y=>nx26440, A0=>
      booth_booth_integrtaion_0_booth_output_21, A1=>nx5134, B0=>nx5114, B1
      =>nx13074);
   ix26444 : nor02ii port map ( Y=>nx26443, A0=>nx5100, A1=>mdr_data_out(21)
   );
   ix5101 : nor02ii port map ( Y=>nx5100, A0=>mdr_data_out(20), A1=>nx5076);
   ix5125 : nor02ii port map ( Y=>nx5124, A0=>mdr_data_out(21), A1=>nx5100);
   ix26454 : xnor2 port map ( Y=>nx26453, A0=>nx5162, A1=>nx13077);
   ix5163 : oai22 port map ( Y=>nx5162, A0=>nx26440, A1=>nx26456, B0=>
      nx26465, B1=>nx35209);
   ix26459 : aoi32 port map ( Y=>nx26458, A0=>nx5144, A1=>nx34681, A2=>
      nx26463, B0=>mdr_data_out(22), B1=>nx34675);
   ix5145 : nand02 port map ( Y=>nx5144, A0=>nx26461, A1=>mdr_data_out(22));
   booth_booth_integrtaion_0_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_22, QB=>nx26465, D=>nx16983, 
      CLK=>clk, R=>rst);
   ix16974 : oai21 port map ( Y=>nx16973, A0=>nx26470, A1=>nx35193, B0=>
      nx26472);
   booth_booth_integrtaion_0_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_23, QB=>nx26470, D=>nx16973, 
      CLK=>clk, R=>rst);
   ix26473 : nand03 port map ( Y=>nx26472, A0=>nx35201, A1=>nx5450, A2=>
      nx35195);
   ix5451 : xnor2 port map ( Y=>nx5450, A0=>nx26475, A1=>nx13079);
   ix26476 : aoi22 port map ( Y=>nx26475, A0=>
      booth_booth_integrtaion_0_booth_output_23, A1=>nx5182, B0=>nx5162, B1
      =>nx13077);
   ix26479 : nor02ii port map ( Y=>nx26478, A0=>nx5148, A1=>mdr_data_out(23)
   );
   ix5149 : nor02ii port map ( Y=>nx5148, A0=>mdr_data_out(22), A1=>nx5124);
   ix5173 : nor02ii port map ( Y=>nx5172, A0=>mdr_data_out(23), A1=>nx5148);
   ix26489 : xnor2 port map ( Y=>nx26488, A0=>nx5210, A1=>nx13081);
   ix5211 : oai22 port map ( Y=>nx5210, A0=>nx26475, A1=>nx26491, B0=>
      nx26500, B1=>nx35211);
   ix26494 : aoi32 port map ( Y=>nx26493, A0=>nx5192, A1=>nx34681, A2=>
      nx26498, B0=>mdr_data_out(24), B1=>nx34675);
   ix5193 : nand02 port map ( Y=>nx5192, A0=>nx26496, A1=>mdr_data_out(24));
   booth_booth_integrtaion_0_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_24, QB=>nx26500, D=>nx16963, 
      CLK=>clk, R=>rst);
   ix16954 : oai21 port map ( Y=>nx16953, A0=>nx26505, A1=>nx35195, B0=>
      nx26507);
   booth_booth_integrtaion_0_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_25, QB=>nx26505, D=>nx16953, 
      CLK=>clk, R=>rst);
   ix26508 : nand03 port map ( Y=>nx26507, A0=>nx35201, A1=>nx5426, A2=>
      nx35195);
   ix5427 : xnor2 port map ( Y=>nx5426, A0=>nx26510, A1=>nx13083);
   ix26511 : aoi22 port map ( Y=>nx26510, A0=>
      booth_booth_integrtaion_0_booth_output_25, A1=>nx5230, B0=>nx5210, B1
      =>nx13081);
   ix26514 : nor02ii port map ( Y=>nx26513, A0=>nx5196, A1=>mdr_data_out(25)
   );
   ix5197 : nor02ii port map ( Y=>nx5196, A0=>mdr_data_out(24), A1=>nx5172);
   ix5221 : nor02ii port map ( Y=>nx5220, A0=>mdr_data_out(25), A1=>nx5196);
   ix26524 : xnor2 port map ( Y=>nx26523, A0=>nx5258, A1=>nx13085);
   ix5259 : oai22 port map ( Y=>nx5258, A0=>nx26510, A1=>nx26526, B0=>
      nx26535, B1=>nx35213);
   ix26529 : aoi32 port map ( Y=>nx26528, A0=>nx5240, A1=>nx34681, A2=>
      nx26533, B0=>mdr_data_out(26), B1=>nx34675);
   ix5241 : nand02 port map ( Y=>nx5240, A0=>nx26531, A1=>mdr_data_out(26));
   booth_booth_integrtaion_0_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_26, QB=>nx26535, D=>nx16943, 
      CLK=>clk, R=>rst);
   ix16934 : oai21 port map ( Y=>nx16933, A0=>nx26540, A1=>nx35195, B0=>
      nx26542);
   booth_booth_integrtaion_0_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_27, QB=>nx26540, D=>nx16933, 
      CLK=>clk, R=>rst);
   ix26543 : nand03 port map ( Y=>nx26542, A0=>nx35201, A1=>nx5402, A2=>
      nx35195);
   ix5403 : xnor2 port map ( Y=>nx5402, A0=>nx26545, A1=>nx13087);
   ix26546 : aoi22 port map ( Y=>nx26545, A0=>
      booth_booth_integrtaion_0_booth_output_27, A1=>nx5278, B0=>nx5258, B1
      =>nx13085);
   ix26549 : nor02ii port map ( Y=>nx26548, A0=>nx5244, A1=>mdr_data_out(27)
   );
   ix5245 : nor02ii port map ( Y=>nx5244, A0=>mdr_data_out(26), A1=>nx5220);
   ix5269 : nor02ii port map ( Y=>nx5268, A0=>mdr_data_out(27), A1=>nx5244);
   ix26559 : xnor2 port map ( Y=>nx26558, A0=>nx5306, A1=>nx13089);
   ix5307 : oai22 port map ( Y=>nx5306, A0=>nx26545, A1=>nx26561, B0=>
      nx26570, B1=>nx35215);
   ix26564 : aoi32 port map ( Y=>nx26563, A0=>nx5288, A1=>nx34681, A2=>
      nx26568, B0=>mdr_data_out(28), B1=>nx34675);
   ix5289 : nand02 port map ( Y=>nx5288, A0=>nx26566, A1=>mdr_data_out(28));
   booth_booth_integrtaion_0_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_28, QB=>nx26570, D=>nx16923, 
      CLK=>clk, R=>rst);
   ix16914 : oai21 port map ( Y=>nx16913, A0=>nx26575, A1=>nx35195, B0=>
      nx26577);
   booth_booth_integrtaion_0_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_29, QB=>nx26575, D=>nx16913, 
      CLK=>clk, R=>rst);
   ix26578 : nand03 port map ( Y=>nx26577, A0=>nx36011, A1=>nx5378, A2=>
      nx35195);
   ix5379 : xnor2 port map ( Y=>nx5378, A0=>nx26580, A1=>nx13090);
   ix26581 : aoi22 port map ( Y=>nx26580, A0=>
      booth_booth_integrtaion_0_booth_output_29, A1=>nx5326, B0=>nx5306, B1
      =>nx13089);
   ix26584 : nor02ii port map ( Y=>nx26583, A0=>nx5292, A1=>mdr_data_out(29)
   );
   ix5293 : nor02ii port map ( Y=>nx5292, A0=>mdr_data_out(28), A1=>nx5268);
   ix5317 : nor02ii port map ( Y=>nx5316, A0=>mdr_data_out(29), A1=>nx5292);
   ix26594 : xnor2 port map ( Y=>nx26593, A0=>nx5354, A1=>nx5364);
   ix5355 : oai22 port map ( Y=>nx5354, A0=>nx26580, A1=>nx26596, B0=>
      nx26605, B1=>nx35217);
   ix26599 : aoi32 port map ( Y=>nx26598, A0=>nx5336, A1=>nx34683, A2=>
      nx26603, B0=>mdr_data_out(30), B1=>nx34677);
   ix5337 : nand02 port map ( Y=>nx5336, A0=>nx26601, A1=>mdr_data_out(30));
   booth_booth_integrtaion_0_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_31, QB=>nx26605, D=>nx16903, 
      CLK=>clk, R=>rst);
   ix26609 : aoi22 port map ( Y=>nx26608, A0=>mdr_data_out(31), A1=>nx34677, 
      B0=>nx34683, B1=>nx5356);
   ix5357 : xnor2 port map ( Y=>nx5356, A0=>mdr_data_out(31), A1=>nx5340);
   ix5341 : nor02ii port map ( Y=>nx5340, A0=>mdr_data_out(30), A1=>nx5316);
   ix26613 : aoi32 port map ( Y=>nx26612, A0=>nx5312, A1=>nx34683, A2=>
      nx26601, B0=>mdr_data_out(29), B1=>nx34677);
   ix26616 : aoi32 port map ( Y=>nx26615, A0=>nx5264, A1=>nx34683, A2=>
      nx26566, B0=>mdr_data_out(27), B1=>nx34677);
   ix26619 : aoi32 port map ( Y=>nx26618, A0=>nx5216, A1=>nx34683, A2=>
      nx26531, B0=>mdr_data_out(25), B1=>nx34677);
   ix26622 : aoi32 port map ( Y=>nx26621, A0=>nx5168, A1=>nx34683, A2=>
      nx26496, B0=>mdr_data_out(23), B1=>nx34677);
   ix26625 : aoi32 port map ( Y=>nx26624, A0=>nx5120, A1=>nx34683, A2=>
      nx26461, B0=>mdr_data_out(21), B1=>nx34677);
   ix26628 : aoi32 port map ( Y=>nx26627, A0=>nx5072, A1=>nx5008, A2=>
      nx26426, B0=>mdr_data_out(19), B1=>nx34679);
   ix26631 : aoi32 port map ( Y=>nx26630, A0=>nx5022, A1=>nx5008, A2=>
      nx26375, B0=>mdr_data_out(17), B1=>nx34679);
   booth_booth_integrtaion_0_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_0_booth_output_16, QB=>nx26356, D=>nx17043, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_0_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_0_15, QB=>nx26634, D=>nx17053, CLK=>clk, 
      R=>rst);
   ix5747 : aoi21 port map ( Y=>nx5746, A0=>label_1_output(0), A1=>nx35731, 
      B0=>nx36387);
   reg_sel_dst_0 : dffr port map ( Q=>sel_dst_0, QB=>OPEN, D=>nx14113, CLK=>
      clk, R=>rst);
   ix14114 : mux21_ni port map ( Y=>nx14113, A0=>sel_dst_0, A1=>nx36201, S0
      =>nx878);
   ix879 : nor03_2x port map ( Y=>nx878, A0=>nx12895, A1=>nx56, A2=>nx26661
   );
   ix26662 : oai21 port map ( Y=>nx26661, A0=>nx25944, A1=>nx35099, B0=>
      nx868);
   ix869 : oai21 port map ( Y=>nx868, A0=>nx26664, A1=>nx26666, B0=>nx172);
   max_calc_reg_ans1_0 : dff port map ( Q=>max_calc_ans1_0, QB=>OPEN, D=>
      nx17583, CLK=>clk);
   ix26676 : nand04 port map ( Y=>nx26675, A0=>nx25940, A1=>max_calc_start, 
      A2=>nx26188, A3=>nx6368);
   ix6369 : aoi21 port map ( Y=>nx6368, A0=>nx35977, A1=>nx36389, B0=>
      max_calc_state_3);
   max_calc_reg_ans6_0 : dff port map ( Q=>max_calc_ans6_0, QB=>OPEN, D=>
      nx17593, CLK=>clk);
   max_calc_reg_ans5_0 : dff port map ( Q=>max_calc_ans5_0, QB=>OPEN, D=>
      nx19623, CLK=>clk);
   ix18154 : oai21 port map ( Y=>nx18153, A0=>nx26693, A1=>nx34747, B0=>
      nx26696);
   max_calc_reg_comparator_fifth_inp1_0 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_0, QB=>nx26693, D=>nx18153, CLK=>clk);
   ix26697 : nand03 port map ( Y=>nx26696, A0=>label_9_output(0), A1=>
      nx34737, A2=>nx34747);
   labelsregfile_label9_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_9_output(0), QB=>OPEN, D=>nx18143, CLK=>clk, R=>rst);
   lat_label_9_input_0 : latch port map ( Q=>label_9_input_0, D=>nx7260, CLK
      =>nx34511);
   ix7261 : oai21 port map ( Y=>nx7260, A0=>nx26702, A1=>nx34409, B0=>
      nx26706);
   reg_label_9_input_state_machine_0 : dffr port map ( Q=>
      label_9_input_state_machine_0, QB=>nx26702, D=>nx18133, CLK=>clk, R=>
      rst);
   ix26707 : oai21 port map ( Y=>nx26706, A0=>nx35755, A1=>label_9_output(0), 
      B0=>nx7248);
   booth_booth_integrtaion_8_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_1, QB=>OPEN, D=>nx18113, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_2, QB=>nx27127, D=>nx18103, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_3, QB=>OPEN, D=>nx18093, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_4, QB=>nx27125, D=>nx18083, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_5, QB=>OPEN, D=>nx18073, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_6, QB=>nx27123, D=>nx18063, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_7, QB=>OPEN, D=>nx18053, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_8, QB=>nx27121, D=>nx18043, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_9, QB=>OPEN, D=>nx18033, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_10, QB=>nx27119, D=>nx18023, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_11, QB=>OPEN, D=>nx18013, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_12, QB=>nx27117, D=>nx18003, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_13, QB=>OPEN, D=>nx17993, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_14, QB=>nx27115, D=>nx17983, CLK=>clk, 
      R=>rst);
   ix26756 : aoi22 port map ( Y=>nx26755, A0=>mdr_data_out(15), A1=>nx34847, 
      B0=>nx7044, B1=>nx7050);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_reg_output_0, QB=>OPEN, 
      D=>nx17623, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_0, QB=>OPEN, D=>nx17609, CLK
      =>clk, S=>nx34467);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_reg_output_9, QB=>OPEN, 
      D=>nx17803, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_9, QB=>OPEN, D=>nx17793, CLK
      =>clk, R=>nx34467);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_8, QB=>OPEN, 
      D=>nx17783, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_8, QB=>OPEN, D=>nx17773, CLK
      =>clk, R=>nx34467);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_7, QB=>OPEN, 
      D=>nx17763, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_7, QB=>OPEN, D=>nx17753, CLK
      =>clk, R=>nx34467);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_6, QB=>OPEN, 
      D=>nx17743, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_6, QB=>OPEN, D=>nx17733, CLK
      =>clk, R=>nx34467);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_5, QB=>OPEN, 
      D=>nx17723, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_5, QB=>OPEN, D=>nx17713, CLK
      =>clk, R=>nx34467);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_4, QB=>OPEN, 
      D=>nx17703, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_4, QB=>OPEN, D=>nx17693, CLK
      =>clk, R=>nx34467);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_3, QB=>OPEN, 
      D=>nx17683, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_3, QB=>OPEN, D=>nx17673, CLK
      =>clk, R=>nx34465);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_2, QB=>OPEN, 
      D=>nx17663, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_2, QB=>OPEN, D=>nx17653, CLK
      =>clk, R=>nx34465);
   booth_booth_integrtaion_8_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_8_shift_Reg_output_1, QB=>OPEN, 
      D=>nx17643, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_8_shift_Reg_count_1, QB=>OPEN, D=>nx17633, CLK
      =>clk, R=>nx34465);
   ix17604 : nand02 port map ( Y=>nx17603, A0=>nx35807, A1=>nx34833);
   booth_booth_integrtaion_8_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx26802, D=>nx17603, CLK=>clk, S=>nx34465);
   ix7045 : nand02 port map ( Y=>nx7044, A0=>nx26823, A1=>nx26835);
   ix26824 : oai21 port map ( Y=>nx26823, A0=>nx34861, A1=>nx34855, B0=>
      mdr_data_out(144));
   ix17814 : oai21 port map ( Y=>nx17813, A0=>nx26828, A1=>nx35301, B0=>
      nx26830);
   booth_booth_integrtaion_8_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx26828, D=>nx17813, CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx26832, D=>nx18123, CLK=>clk, R=>rst);
   ix26840 : xnor2 port map ( Y=>nx26839, A0=>nx6514, A1=>nx13123);
   ix17954 : oai21 port map ( Y=>nx17953, A0=>nx26845, A1=>nx35301, B0=>
      nx26847);
   booth_booth_integrtaion_8_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_17, QB=>nx26845, D=>nx17953, 
      CLK=>clk, R=>rst);
   ix26848 : nand03 port map ( Y=>nx26847, A0=>nx35309, A1=>nx7022, A2=>
      nx36031);
   ix7023 : xnor2 port map ( Y=>nx7022, A0=>nx26850, A1=>nx13125);
   ix26851 : aoi22 port map ( Y=>nx26850, A0=>
      booth_booth_integrtaion_8_booth_output_17, A1=>nx6538, B0=>nx6514, B1
      =>nx13123);
   ix6523 : nand02 port map ( Y=>nx6522, A0=>mdr_data_out(145), A1=>
      mdr_data_out(144));
   ix26855 : or02 port map ( Y=>nx26854, A0=>mdr_data_out(144), A1=>
      mdr_data_out(145));
   ix26861 : xnor2 port map ( Y=>nx26860, A0=>nx6566, A1=>nx13127);
   ix6567 : oai22 port map ( Y=>nx6566, A0=>nx26850, A1=>nx26863, B0=>
      nx26870, B1=>nx35313);
   ix26866 : aoi32 port map ( Y=>nx26865, A0=>nx6548, A1=>nx34861, A2=>
      nx26868, B0=>mdr_data_out(146), B1=>nx34855);
   ix6549 : oai21 port map ( Y=>nx6548, A0=>mdr_data_out(144), A1=>
      mdr_data_out(145), B0=>mdr_data_out(146));
   booth_booth_integrtaion_8_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_18, QB=>nx26870, D=>nx17943, 
      CLK=>clk, R=>rst);
   ix17934 : oai21 port map ( Y=>nx17933, A0=>nx26875, A1=>nx35301, B0=>
      nx26877);
   booth_booth_integrtaion_8_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_19, QB=>nx26875, D=>nx17933, 
      CLK=>clk, R=>rst);
   ix26878 : nand03 port map ( Y=>nx26877, A0=>nx35309, A1=>nx6998, A2=>
      nx36031);
   ix6999 : xnor2 port map ( Y=>nx6998, A0=>nx26880, A1=>nx13129);
   ix26881 : aoi22 port map ( Y=>nx26880, A0=>
      booth_booth_integrtaion_8_booth_output_19, A1=>nx6586, B0=>nx6566, B1
      =>nx13127);
   ix26884 : nor02ii port map ( Y=>nx26883, A0=>nx6552, A1=>
      mdr_data_out(147));
   ix6553 : nor03_2x port map ( Y=>nx6552, A0=>mdr_data_out(146), A1=>
      mdr_data_out(144), A2=>mdr_data_out(145));
   ix6577 : nor04 port map ( Y=>nx6576, A0=>mdr_data_out(147), A1=>
      mdr_data_out(146), A2=>mdr_data_out(144), A3=>mdr_data_out(145));
   ix26898 : xnor2 port map ( Y=>nx26897, A0=>nx6614, A1=>nx13131);
   ix6615 : oai22 port map ( Y=>nx6614, A0=>nx26880, A1=>nx26900, B0=>
      nx26909, B1=>nx35315);
   ix26903 : aoi32 port map ( Y=>nx26902, A0=>nx6596, A1=>nx34861, A2=>
      nx26907, B0=>mdr_data_out(148), B1=>nx34855);
   ix6597 : nand02 port map ( Y=>nx6596, A0=>nx26905, A1=>mdr_data_out(148)
   );
   booth_booth_integrtaion_8_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_20, QB=>nx26909, D=>nx17923, 
      CLK=>clk, R=>rst);
   ix17914 : oai21 port map ( Y=>nx17913, A0=>nx26914, A1=>nx35301, B0=>
      nx26916);
   booth_booth_integrtaion_8_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_21, QB=>nx26914, D=>nx17913, 
      CLK=>clk, R=>rst);
   ix26917 : nand03 port map ( Y=>nx26916, A0=>nx35309, A1=>nx6974, A2=>
      nx36031);
   ix6975 : xnor2 port map ( Y=>nx6974, A0=>nx26919, A1=>nx13133);
   ix26920 : aoi22 port map ( Y=>nx26919, A0=>
      booth_booth_integrtaion_8_booth_output_21, A1=>nx6634, B0=>nx6614, B1
      =>nx13131);
   ix26923 : nor02ii port map ( Y=>nx26922, A0=>nx6600, A1=>
      mdr_data_out(149));
   ix6601 : nor02ii port map ( Y=>nx6600, A0=>mdr_data_out(148), A1=>nx6576
   );
   ix6625 : nor02ii port map ( Y=>nx6624, A0=>mdr_data_out(149), A1=>nx6600
   );
   ix26933 : xnor2 port map ( Y=>nx26932, A0=>nx6662, A1=>nx13135);
   ix6663 : oai22 port map ( Y=>nx6662, A0=>nx26919, A1=>nx26935, B0=>
      nx26944, B1=>nx35317);
   ix26938 : aoi32 port map ( Y=>nx26937, A0=>nx6644, A1=>nx34861, A2=>
      nx26942, B0=>mdr_data_out(150), B1=>nx34855);
   ix6645 : nand02 port map ( Y=>nx6644, A0=>nx26940, A1=>mdr_data_out(150)
   );
   booth_booth_integrtaion_8_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_22, QB=>nx26944, D=>nx17903, 
      CLK=>clk, R=>rst);
   ix17894 : oai21 port map ( Y=>nx17893, A0=>nx26949, A1=>nx35301, B0=>
      nx26951);
   booth_booth_integrtaion_8_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_23, QB=>nx26949, D=>nx17893, 
      CLK=>clk, R=>rst);
   ix26952 : nand03 port map ( Y=>nx26951, A0=>nx35309, A1=>nx6950, A2=>
      nx35303);
   ix6951 : xnor2 port map ( Y=>nx6950, A0=>nx26954, A1=>nx13137);
   ix26955 : aoi22 port map ( Y=>nx26954, A0=>
      booth_booth_integrtaion_8_booth_output_23, A1=>nx6682, B0=>nx6662, B1
      =>nx13135);
   ix26958 : nor02ii port map ( Y=>nx26957, A0=>nx6648, A1=>
      mdr_data_out(151));
   ix6649 : nor02ii port map ( Y=>nx6648, A0=>mdr_data_out(150), A1=>nx6624
   );
   ix6673 : nor02ii port map ( Y=>nx6672, A0=>mdr_data_out(151), A1=>nx6648
   );
   ix26968 : xnor2 port map ( Y=>nx26967, A0=>nx6710, A1=>nx13138);
   ix6711 : oai22 port map ( Y=>nx6710, A0=>nx26954, A1=>nx26970, B0=>
      nx26979, B1=>nx35319);
   ix26973 : aoi32 port map ( Y=>nx26972, A0=>nx6692, A1=>nx34861, A2=>
      nx26977, B0=>mdr_data_out(152), B1=>nx34855);
   ix6693 : nand02 port map ( Y=>nx6692, A0=>nx26975, A1=>mdr_data_out(152)
   );
   booth_booth_integrtaion_8_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_24, QB=>nx26979, D=>nx17883, 
      CLK=>clk, R=>rst);
   ix17874 : oai21 port map ( Y=>nx17873, A0=>nx26984, A1=>nx35303, B0=>
      nx26986);
   booth_booth_integrtaion_8_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_25, QB=>nx26984, D=>nx17873, 
      CLK=>clk, R=>rst);
   ix26987 : nand03 port map ( Y=>nx26986, A0=>nx35309, A1=>nx6926, A2=>
      nx35303);
   ix6927 : xnor2 port map ( Y=>nx6926, A0=>nx26989, A1=>nx13139);
   ix26990 : aoi22 port map ( Y=>nx26989, A0=>
      booth_booth_integrtaion_8_booth_output_25, A1=>nx6730, B0=>nx6710, B1
      =>nx13138);
   ix26993 : nor02ii port map ( Y=>nx26992, A0=>nx6696, A1=>
      mdr_data_out(153));
   ix6697 : nor02ii port map ( Y=>nx6696, A0=>mdr_data_out(152), A1=>nx6672
   );
   ix6721 : nor02ii port map ( Y=>nx6720, A0=>mdr_data_out(153), A1=>nx6696
   );
   ix27003 : xnor2 port map ( Y=>nx27002, A0=>nx6758, A1=>nx13141);
   ix6759 : oai22 port map ( Y=>nx6758, A0=>nx26989, A1=>nx27005, B0=>
      nx27014, B1=>nx35321);
   ix27008 : aoi32 port map ( Y=>nx27007, A0=>nx6740, A1=>nx34861, A2=>
      nx27012, B0=>mdr_data_out(154), B1=>nx34855);
   ix6741 : nand02 port map ( Y=>nx6740, A0=>nx27010, A1=>mdr_data_out(154)
   );
   booth_booth_integrtaion_8_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_26, QB=>nx27014, D=>nx17863, 
      CLK=>clk, R=>rst);
   ix17854 : oai21 port map ( Y=>nx17853, A0=>nx27019, A1=>nx35303, B0=>
      nx27021);
   booth_booth_integrtaion_8_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_27, QB=>nx27019, D=>nx17853, 
      CLK=>clk, R=>rst);
   ix27022 : nand03 port map ( Y=>nx27021, A0=>nx35309, A1=>nx6902, A2=>
      nx35303);
   ix6903 : xnor2 port map ( Y=>nx6902, A0=>nx27024, A1=>nx13143);
   ix27025 : aoi22 port map ( Y=>nx27024, A0=>
      booth_booth_integrtaion_8_booth_output_27, A1=>nx6778, B0=>nx6758, B1
      =>nx13141);
   ix27028 : nor02ii port map ( Y=>nx27027, A0=>nx6744, A1=>
      mdr_data_out(155));
   ix6745 : nor02ii port map ( Y=>nx6744, A0=>mdr_data_out(154), A1=>nx6720
   );
   ix6769 : nor02ii port map ( Y=>nx6768, A0=>mdr_data_out(155), A1=>nx6744
   );
   ix27038 : xnor2 port map ( Y=>nx27037, A0=>nx6806, A1=>nx13145);
   ix6807 : oai22 port map ( Y=>nx6806, A0=>nx27024, A1=>nx27040, B0=>
      nx27049, B1=>nx35323);
   ix27043 : aoi32 port map ( Y=>nx27042, A0=>nx6788, A1=>nx34861, A2=>
      nx27047, B0=>mdr_data_out(156), B1=>nx34855);
   ix6789 : nand02 port map ( Y=>nx6788, A0=>nx27045, A1=>mdr_data_out(156)
   );
   booth_booth_integrtaion_8_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_28, QB=>nx27049, D=>nx17843, 
      CLK=>clk, R=>rst);
   ix17834 : oai21 port map ( Y=>nx17833, A0=>nx27054, A1=>nx35303, B0=>
      nx27056);
   booth_booth_integrtaion_8_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_29, QB=>nx27054, D=>nx17833, 
      CLK=>clk, R=>rst);
   ix27057 : nand03 port map ( Y=>nx27056, A0=>nx36039, A1=>nx6878, A2=>
      nx35303);
   ix6879 : xnor2 port map ( Y=>nx6878, A0=>nx27059, A1=>nx13146);
   ix27060 : aoi22 port map ( Y=>nx27059, A0=>
      booth_booth_integrtaion_8_booth_output_29, A1=>nx6826, B0=>nx6806, B1
      =>nx13145);
   ix27063 : nor02ii port map ( Y=>nx27062, A0=>nx6792, A1=>
      mdr_data_out(157));
   ix6793 : nor02ii port map ( Y=>nx6792, A0=>mdr_data_out(156), A1=>nx6768
   );
   ix6817 : nor02ii port map ( Y=>nx6816, A0=>mdr_data_out(157), A1=>nx6792
   );
   ix27073 : xnor2 port map ( Y=>nx27072, A0=>nx6854, A1=>nx6864);
   ix6855 : oai22 port map ( Y=>nx6854, A0=>nx27059, A1=>nx27075, B0=>
      nx27084, B1=>nx35325);
   ix27078 : aoi32 port map ( Y=>nx27077, A0=>nx6836, A1=>nx34863, A2=>
      nx27082, B0=>mdr_data_out(158), B1=>nx34857);
   ix6837 : nand02 port map ( Y=>nx6836, A0=>nx27080, A1=>mdr_data_out(158)
   );
   booth_booth_integrtaion_8_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_31, QB=>nx27084, D=>nx17823, 
      CLK=>clk, R=>rst);
   ix27088 : aoi22 port map ( Y=>nx27087, A0=>mdr_data_out(159), A1=>nx34857, 
      B0=>nx34863, B1=>nx6856);
   ix6857 : xnor2 port map ( Y=>nx6856, A0=>mdr_data_out(159), A1=>nx6840);
   ix6841 : nor02ii port map ( Y=>nx6840, A0=>mdr_data_out(158), A1=>nx6816
   );
   ix27092 : aoi32 port map ( Y=>nx27091, A0=>nx6812, A1=>nx34863, A2=>
      nx27080, B0=>mdr_data_out(157), B1=>nx34857);
   ix27095 : aoi32 port map ( Y=>nx27094, A0=>nx6764, A1=>nx34863, A2=>
      nx27045, B0=>mdr_data_out(155), B1=>nx34857);
   ix27098 : aoi32 port map ( Y=>nx27097, A0=>nx6716, A1=>nx34863, A2=>
      nx27010, B0=>mdr_data_out(153), B1=>nx34857);
   ix27101 : aoi32 port map ( Y=>nx27100, A0=>nx6668, A1=>nx34863, A2=>
      nx26975, B0=>mdr_data_out(151), B1=>nx34857);
   ix27104 : aoi32 port map ( Y=>nx27103, A0=>nx6620, A1=>nx34863, A2=>
      nx26940, B0=>mdr_data_out(149), B1=>nx34857);
   ix27107 : aoi32 port map ( Y=>nx27106, A0=>nx6572, A1=>nx6508, A2=>
      nx26905, B0=>mdr_data_out(147), B1=>nx34859);
   ix27110 : aoi32 port map ( Y=>nx27109, A0=>nx6522, A1=>nx6508, A2=>
      nx26854, B0=>mdr_data_out(145), B1=>nx34859);
   booth_booth_integrtaion_8_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_8_booth_output_16, QB=>nx26835, D=>nx17963, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_8_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_8_15, QB=>nx27113, D=>nx17973, CLK=>clk, 
      R=>rst);
   ix7249 : aoi21 port map ( Y=>nx7248, A0=>label_9_output(0), A1=>nx35755, 
      B0=>nx36387);
   ix19554 : oai21 port map ( Y=>nx19553, A0=>nx27133, A1=>nx34747, B0=>
      nx27135);
   max_calc_reg_comparator_fifth_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx27133, D=>nx19553, CLK=>clk);
   ix27136 : nand03 port map ( Y=>nx27135, A0=>label_10_output(0), A1=>
      nx34737, A2=>nx34747);
   labelsregfile_label10_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_10_output(0), QB=>OPEN, D=>nx18713, CLK=>clk, R=>rst);
   lat_label_10_input_0 : latch port map ( Q=>label_10_input_0, D=>nx8138, 
      CLK=>nx34511);
   ix8139 : oai21 port map ( Y=>nx8138, A0=>nx27141, A1=>nx34409, B0=>
      nx27145);
   reg_label_10_input_state_machine_0 : dffr port map ( Q=>
      label_10_input_state_machine_0, QB=>nx27141, D=>nx18703, CLK=>clk, R=>
      rst);
   ix27146 : oai21 port map ( Y=>nx27145, A0=>nx35759, A1=>
      label_10_output(0), B0=>nx8126);
   booth_booth_integrtaion_9_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_1, QB=>OPEN, D=>nx18683, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_2, QB=>nx27566, D=>nx18673, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_3, QB=>OPEN, D=>nx18663, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_4, QB=>nx27564, D=>nx18653, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_5, QB=>OPEN, D=>nx18643, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_6, QB=>nx27562, D=>nx18633, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_7, QB=>OPEN, D=>nx18623, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_8, QB=>nx27560, D=>nx18613, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_9, QB=>OPEN, D=>nx18603, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_10, QB=>nx27558, D=>nx18593, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_11, QB=>OPEN, D=>nx18583, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_12, QB=>nx27556, D=>nx18573, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_13, QB=>OPEN, D=>nx18563, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_14, QB=>nx27554, D=>nx18553, CLK=>clk, 
      R=>rst);
   ix27195 : aoi22 port map ( Y=>nx27194, A0=>mdr_data_out(15), A1=>nx34879, 
      B0=>nx7924, B1=>nx7930);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_reg_output_0, QB=>OPEN, 
      D=>nx18193, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_0, QB=>OPEN, D=>nx18179, CLK
      =>clk, S=>nx34471);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_reg_output_9, QB=>OPEN, 
      D=>nx18373, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_9, QB=>OPEN, D=>nx18363, CLK
      =>clk, R=>nx34471);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_8, QB=>OPEN, 
      D=>nx18353, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_8, QB=>OPEN, D=>nx18343, CLK
      =>clk, R=>nx34471);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_7, QB=>OPEN, 
      D=>nx18333, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_7, QB=>OPEN, D=>nx18323, CLK
      =>clk, R=>nx34471);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_6, QB=>OPEN, 
      D=>nx18313, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_6, QB=>OPEN, D=>nx18303, CLK
      =>clk, R=>nx34469);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_5, QB=>OPEN, 
      D=>nx18293, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_5, QB=>OPEN, D=>nx18283, CLK
      =>clk, R=>nx34469);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_4, QB=>OPEN, 
      D=>nx18273, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_4, QB=>OPEN, D=>nx18263, CLK
      =>clk, R=>nx34469);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_3, QB=>OPEN, 
      D=>nx18253, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_3, QB=>OPEN, D=>nx18243, CLK
      =>clk, R=>nx34469);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_2, QB=>OPEN, 
      D=>nx18233, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_2, QB=>OPEN, D=>nx18223, CLK
      =>clk, R=>nx34469);
   booth_booth_integrtaion_9_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_9_shift_Reg_output_1, QB=>OPEN, 
      D=>nx18213, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_9_shift_Reg_count_1, QB=>OPEN, D=>nx18203, CLK
      =>clk, R=>nx34469);
   ix18174 : nand02 port map ( Y=>nx18173, A0=>nx35811, A1=>nx34865);
   booth_booth_integrtaion_9_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx27241, D=>nx18173, CLK=>clk, S=>nx34469);
   ix7925 : nand02 port map ( Y=>nx7924, A0=>nx27262, A1=>nx27274);
   ix27263 : oai21 port map ( Y=>nx27262, A0=>nx34893, A1=>nx34887, B0=>
      mdr_data_out(160));
   ix18384 : oai21 port map ( Y=>nx18383, A0=>nx27267, A1=>nx35327, B0=>
      nx27269);
   booth_booth_integrtaion_9_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx27267, D=>nx18383, CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx27271, D=>nx18693, CLK=>clk, R=>rst);
   ix27279 : xnor2 port map ( Y=>nx27278, A0=>nx7394, A1=>nx13149);
   ix18524 : oai21 port map ( Y=>nx18523, A0=>nx27284, A1=>nx35327, B0=>
      nx27286);
   booth_booth_integrtaion_9_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_17, QB=>nx27284, D=>nx18523, 
      CLK=>clk, R=>rst);
   ix27287 : nand03 port map ( Y=>nx27286, A0=>nx35335, A1=>nx7902, A2=>
      nx36047);
   ix7903 : xnor2 port map ( Y=>nx7902, A0=>nx27289, A1=>nx13151);
   ix27290 : aoi22 port map ( Y=>nx27289, A0=>
      booth_booth_integrtaion_9_booth_output_17, A1=>nx7418, B0=>nx7394, B1
      =>nx13149);
   ix7403 : nand02 port map ( Y=>nx7402, A0=>mdr_data_out(161), A1=>
      mdr_data_out(160));
   ix27294 : or02 port map ( Y=>nx27293, A0=>mdr_data_out(160), A1=>
      mdr_data_out(161));
   ix27300 : xnor2 port map ( Y=>nx27299, A0=>nx7446, A1=>nx13153);
   ix7447 : oai22 port map ( Y=>nx7446, A0=>nx27289, A1=>nx27302, B0=>
      nx27309, B1=>nx35339);
   ix27305 : aoi32 port map ( Y=>nx27304, A0=>nx7428, A1=>nx34893, A2=>
      nx27307, B0=>mdr_data_out(162), B1=>nx34887);
   ix7429 : oai21 port map ( Y=>nx7428, A0=>mdr_data_out(160), A1=>
      mdr_data_out(161), B0=>mdr_data_out(162));
   booth_booth_integrtaion_9_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_18, QB=>nx27309, D=>nx18513, 
      CLK=>clk, R=>rst);
   ix18504 : oai21 port map ( Y=>nx18503, A0=>nx27314, A1=>nx35327, B0=>
      nx27316);
   booth_booth_integrtaion_9_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_19, QB=>nx27314, D=>nx18503, 
      CLK=>clk, R=>rst);
   ix27317 : nand03 port map ( Y=>nx27316, A0=>nx35335, A1=>nx7878, A2=>
      nx36047);
   ix7879 : xnor2 port map ( Y=>nx7878, A0=>nx27319, A1=>nx13155);
   ix27320 : aoi22 port map ( Y=>nx27319, A0=>
      booth_booth_integrtaion_9_booth_output_19, A1=>nx7466, B0=>nx7446, B1
      =>nx13153);
   ix27323 : nor02ii port map ( Y=>nx27322, A0=>nx7432, A1=>
      mdr_data_out(163));
   ix7433 : nor03_2x port map ( Y=>nx7432, A0=>mdr_data_out(162), A1=>
      mdr_data_out(160), A2=>mdr_data_out(161));
   ix7457 : nor04 port map ( Y=>nx7456, A0=>mdr_data_out(163), A1=>
      mdr_data_out(162), A2=>mdr_data_out(160), A3=>mdr_data_out(161));
   ix27337 : xnor2 port map ( Y=>nx27336, A0=>nx7494, A1=>nx13157);
   ix7495 : oai22 port map ( Y=>nx7494, A0=>nx27319, A1=>nx27339, B0=>
      nx27348, B1=>nx35341);
   ix27342 : aoi32 port map ( Y=>nx27341, A0=>nx7476, A1=>nx34893, A2=>
      nx27346, B0=>mdr_data_out(164), B1=>nx34887);
   ix7477 : nand02 port map ( Y=>nx7476, A0=>nx27344, A1=>mdr_data_out(164)
   );
   booth_booth_integrtaion_9_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_20, QB=>nx27348, D=>nx18493, 
      CLK=>clk, R=>rst);
   ix18484 : oai21 port map ( Y=>nx18483, A0=>nx27353, A1=>nx35327, B0=>
      nx27355);
   booth_booth_integrtaion_9_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_21, QB=>nx27353, D=>nx18483, 
      CLK=>clk, R=>rst);
   ix27356 : nand03 port map ( Y=>nx27355, A0=>nx35335, A1=>nx7854, A2=>
      nx36047);
   ix7855 : xnor2 port map ( Y=>nx7854, A0=>nx27358, A1=>nx13159);
   ix27359 : aoi22 port map ( Y=>nx27358, A0=>
      booth_booth_integrtaion_9_booth_output_21, A1=>nx7514, B0=>nx7494, B1
      =>nx13157);
   ix27362 : nor02ii port map ( Y=>nx27361, A0=>nx7480, A1=>
      mdr_data_out(165));
   ix7481 : nor02ii port map ( Y=>nx7480, A0=>mdr_data_out(164), A1=>nx7456
   );
   ix7505 : nor02ii port map ( Y=>nx7504, A0=>mdr_data_out(165), A1=>nx7480
   );
   ix27372 : xnor2 port map ( Y=>nx27371, A0=>nx7542, A1=>nx13161);
   ix7543 : oai22 port map ( Y=>nx7542, A0=>nx27358, A1=>nx27374, B0=>
      nx27383, B1=>nx35343);
   ix27377 : aoi32 port map ( Y=>nx27376, A0=>nx7524, A1=>nx34893, A2=>
      nx27381, B0=>mdr_data_out(166), B1=>nx34887);
   ix7525 : nand02 port map ( Y=>nx7524, A0=>nx27379, A1=>mdr_data_out(166)
   );
   booth_booth_integrtaion_9_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_22, QB=>nx27383, D=>nx18473, 
      CLK=>clk, R=>rst);
   ix18464 : oai21 port map ( Y=>nx18463, A0=>nx27388, A1=>nx35327, B0=>
      nx27390);
   booth_booth_integrtaion_9_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_23, QB=>nx27388, D=>nx18463, 
      CLK=>clk, R=>rst);
   ix27391 : nand03 port map ( Y=>nx27390, A0=>nx35335, A1=>nx7830, A2=>
      nx35329);
   ix7831 : xnor2 port map ( Y=>nx7830, A0=>nx27393, A1=>nx13162);
   ix27394 : aoi22 port map ( Y=>nx27393, A0=>
      booth_booth_integrtaion_9_booth_output_23, A1=>nx7562, B0=>nx7542, B1
      =>nx13161);
   ix27397 : nor02ii port map ( Y=>nx27396, A0=>nx7528, A1=>
      mdr_data_out(167));
   ix7529 : nor02ii port map ( Y=>nx7528, A0=>mdr_data_out(166), A1=>nx7504
   );
   ix7553 : nor02ii port map ( Y=>nx7552, A0=>mdr_data_out(167), A1=>nx7528
   );
   ix27407 : xnor2 port map ( Y=>nx27406, A0=>nx7590, A1=>nx13163);
   ix7591 : oai22 port map ( Y=>nx7590, A0=>nx27393, A1=>nx27409, B0=>
      nx27418, B1=>nx35345);
   ix27412 : aoi32 port map ( Y=>nx27411, A0=>nx7572, A1=>nx34893, A2=>
      nx27416, B0=>mdr_data_out(168), B1=>nx34887);
   ix7573 : nand02 port map ( Y=>nx7572, A0=>nx27414, A1=>mdr_data_out(168)
   );
   booth_booth_integrtaion_9_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_24, QB=>nx27418, D=>nx18453, 
      CLK=>clk, R=>rst);
   ix18444 : oai21 port map ( Y=>nx18443, A0=>nx27423, A1=>nx35329, B0=>
      nx27425);
   booth_booth_integrtaion_9_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_25, QB=>nx27423, D=>nx18443, 
      CLK=>clk, R=>rst);
   ix27426 : nand03 port map ( Y=>nx27425, A0=>nx35335, A1=>nx7806, A2=>
      nx35329);
   ix7807 : xnor2 port map ( Y=>nx7806, A0=>nx27428, A1=>nx13165);
   ix27429 : aoi22 port map ( Y=>nx27428, A0=>
      booth_booth_integrtaion_9_booth_output_25, A1=>nx7610, B0=>nx7590, B1
      =>nx13163);
   ix27432 : nor02ii port map ( Y=>nx27431, A0=>nx7576, A1=>
      mdr_data_out(169));
   ix7577 : nor02ii port map ( Y=>nx7576, A0=>mdr_data_out(168), A1=>nx7552
   );
   ix7601 : nor02ii port map ( Y=>nx7600, A0=>mdr_data_out(169), A1=>nx7576
   );
   ix27442 : xnor2 port map ( Y=>nx27441, A0=>nx7638, A1=>nx13167);
   ix7639 : oai22 port map ( Y=>nx7638, A0=>nx27428, A1=>nx27444, B0=>
      nx27453, B1=>nx35347);
   ix27447 : aoi32 port map ( Y=>nx27446, A0=>nx7620, A1=>nx34893, A2=>
      nx27451, B0=>mdr_data_out(170), B1=>nx34887);
   ix7621 : nand02 port map ( Y=>nx7620, A0=>nx27449, A1=>mdr_data_out(170)
   );
   booth_booth_integrtaion_9_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_26, QB=>nx27453, D=>nx18433, 
      CLK=>clk, R=>rst);
   ix18424 : oai21 port map ( Y=>nx18423, A0=>nx27458, A1=>nx35329, B0=>
      nx27460);
   booth_booth_integrtaion_9_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_27, QB=>nx27458, D=>nx18423, 
      CLK=>clk, R=>rst);
   ix27461 : nand03 port map ( Y=>nx27460, A0=>nx35335, A1=>nx7782, A2=>
      nx35329);
   ix7783 : xnor2 port map ( Y=>nx7782, A0=>nx27463, A1=>nx13169);
   ix27464 : aoi22 port map ( Y=>nx27463, A0=>
      booth_booth_integrtaion_9_booth_output_27, A1=>nx7658, B0=>nx7638, B1
      =>nx13167);
   ix27467 : nor02ii port map ( Y=>nx27466, A0=>nx7624, A1=>
      mdr_data_out(171));
   ix7625 : nor02ii port map ( Y=>nx7624, A0=>mdr_data_out(170), A1=>nx7600
   );
   ix7649 : nor02ii port map ( Y=>nx7648, A0=>mdr_data_out(171), A1=>nx7624
   );
   ix27477 : xnor2 port map ( Y=>nx27476, A0=>nx7686, A1=>nx13170);
   ix7687 : oai22 port map ( Y=>nx7686, A0=>nx27463, A1=>nx27479, B0=>
      nx27488, B1=>nx35349);
   ix27482 : aoi32 port map ( Y=>nx27481, A0=>nx7668, A1=>nx34893, A2=>
      nx27486, B0=>mdr_data_out(172), B1=>nx34887);
   ix7669 : nand02 port map ( Y=>nx7668, A0=>nx27484, A1=>mdr_data_out(172)
   );
   booth_booth_integrtaion_9_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_28, QB=>nx27488, D=>nx18413, 
      CLK=>clk, R=>rst);
   ix18404 : oai21 port map ( Y=>nx18403, A0=>nx27493, A1=>nx35329, B0=>
      nx27495);
   booth_booth_integrtaion_9_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_29, QB=>nx27493, D=>nx18403, 
      CLK=>clk, R=>rst);
   ix27496 : nand03 port map ( Y=>nx27495, A0=>nx36055, A1=>nx7758, A2=>
      nx35329);
   ix7759 : xnor2 port map ( Y=>nx7758, A0=>nx27498, A1=>nx13171);
   ix27499 : aoi22 port map ( Y=>nx27498, A0=>
      booth_booth_integrtaion_9_booth_output_29, A1=>nx7706, B0=>nx7686, B1
      =>nx13170);
   ix27502 : nor02ii port map ( Y=>nx27501, A0=>nx7672, A1=>
      mdr_data_out(173));
   ix7673 : nor02ii port map ( Y=>nx7672, A0=>mdr_data_out(172), A1=>nx7648
   );
   ix7697 : nor02ii port map ( Y=>nx7696, A0=>mdr_data_out(173), A1=>nx7672
   );
   ix27512 : xnor2 port map ( Y=>nx27511, A0=>nx7734, A1=>nx7744);
   ix7735 : oai22 port map ( Y=>nx7734, A0=>nx27498, A1=>nx27514, B0=>
      nx27523, B1=>nx35351);
   ix27517 : aoi32 port map ( Y=>nx27516, A0=>nx7716, A1=>nx34895, A2=>
      nx27521, B0=>mdr_data_out(174), B1=>nx34889);
   ix7717 : nand02 port map ( Y=>nx7716, A0=>nx27519, A1=>mdr_data_out(174)
   );
   booth_booth_integrtaion_9_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_31, QB=>nx27523, D=>nx18393, 
      CLK=>clk, R=>rst);
   ix27527 : aoi22 port map ( Y=>nx27526, A0=>mdr_data_out(175), A1=>nx34889, 
      B0=>nx34895, B1=>nx7736);
   ix7737 : xnor2 port map ( Y=>nx7736, A0=>mdr_data_out(175), A1=>nx7720);
   ix7721 : nor02ii port map ( Y=>nx7720, A0=>mdr_data_out(174), A1=>nx7696
   );
   ix27531 : aoi32 port map ( Y=>nx27530, A0=>nx7692, A1=>nx34895, A2=>
      nx27519, B0=>mdr_data_out(173), B1=>nx34889);
   ix27534 : aoi32 port map ( Y=>nx27533, A0=>nx7644, A1=>nx34895, A2=>
      nx27484, B0=>mdr_data_out(171), B1=>nx34889);
   ix27537 : aoi32 port map ( Y=>nx27536, A0=>nx7596, A1=>nx34895, A2=>
      nx27449, B0=>mdr_data_out(169), B1=>nx34889);
   ix27540 : aoi32 port map ( Y=>nx27539, A0=>nx7548, A1=>nx34895, A2=>
      nx27414, B0=>mdr_data_out(167), B1=>nx34889);
   ix27543 : aoi32 port map ( Y=>nx27542, A0=>nx7500, A1=>nx34895, A2=>
      nx27379, B0=>mdr_data_out(165), B1=>nx34889);
   ix27546 : aoi32 port map ( Y=>nx27545, A0=>nx7452, A1=>nx7388, A2=>
      nx27344, B0=>mdr_data_out(163), B1=>nx34891);
   ix27549 : aoi32 port map ( Y=>nx27548, A0=>nx7402, A1=>nx7388, A2=>
      nx27293, B0=>mdr_data_out(161), B1=>nx34891);
   booth_booth_integrtaion_9_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_9_booth_output_16, QB=>nx27274, D=>nx18533, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_9_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_9_15, QB=>nx27552, D=>nx18543, CLK=>clk, 
      R=>rst);
   ix8127 : aoi21 port map ( Y=>nx8126, A0=>label_10_output(0), A1=>nx35759, 
      B0=>nx36387);
   ix9491 : xnor2 port map ( Y=>nx9490, A0=>nx27571, A1=>nx9488);
   ix27572 : aoi22 port map ( Y=>nx27571, A0=>nx27573, A1=>
      max_calc_comparator_fifth_inp1_14, B0=>nx9044, B1=>nx9398);
   max_calc_reg_comparator_fifth_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx27573, D=>nx18993, CLK=>clk);
   ix18994 : oai21 port map ( Y=>nx18993, A0=>nx27573, A1=>nx34747, B0=>
      nx27576);
   labelsregfile_label10_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_10_output(14), QB=>nx27760, D=>nx18983, CLK=>clk, R=>rst);
   lat_label_10_input_14 : latch port map ( Q=>label_10_input_14, D=>nx8574, 
      CLK=>nx34515);
   reg_label_10_input_state_machine_14 : dffr port map ( Q=>
      label_10_input_state_machine_14, QB=>OPEN, D=>nx18163, CLK=>clk, R=>
      rst);
   ix8571 : xor2 port map ( Y=>nx8570, A0=>nx27586, A1=>nx27758);
   ix27587 : aoi22 port map ( Y=>nx27586, A0=>label_10_output(13), A1=>
      booth_booth_integration_output_9_13, B0=>nx8534, B1=>nx13199);
   labelsregfile_label10_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_10_output(13), QB=>OPEN, D=>nx18973, CLK=>clk, R=>rst);
   lat_label_10_input_13 : latch port map ( Q=>label_10_input_13, D=>nx8548, 
      CLK=>nx34515);
   reg_label_10_input_state_machine_13 : dffr port map ( Q=>
      label_10_input_state_machine_13, QB=>OPEN, D=>nx18963, CLK=>clk, R=>
      rst);
   ix8545 : xnor2 port map ( Y=>nx8544, A0=>nx8534, A1=>nx27754);
   ix8535 : oai22 port map ( Y=>nx8534, A0=>nx27597, A1=>nx27743, B0=>
      nx27753, B1=>nx27556);
   ix27598 : aoi22 port map ( Y=>nx27597, A0=>label_10_output(11), A1=>
      booth_booth_integration_output_9_11, B0=>nx8470, B1=>nx13195);
   labelsregfile_label10_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_10_output(11), QB=>OPEN, D=>nx18933, CLK=>clk, R=>rst);
   lat_label_10_input_11 : latch port map ( Q=>label_10_input_11, D=>nx8484, 
      CLK=>nx34513);
   reg_label_10_input_state_machine_11 : dffr port map ( Q=>
      label_10_input_state_machine_11, QB=>OPEN, D=>nx18923, CLK=>clk, R=>
      rst);
   ix8481 : xnor2 port map ( Y=>nx8480, A0=>nx8470, A1=>nx27739);
   ix8471 : oai22 port map ( Y=>nx8470, A0=>nx27608, A1=>nx27728, B0=>
      nx27738, B1=>nx27558);
   ix27609 : aoi22 port map ( Y=>nx27608, A0=>label_10_output(9), A1=>
      booth_booth_integration_output_9_9, B0=>nx8406, B1=>nx13191);
   labelsregfile_label10_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_10_output(9), QB=>OPEN, D=>nx18893, CLK=>clk, R=>rst);
   lat_label_10_input_9 : latch port map ( Q=>label_10_input_9, D=>nx8420, 
      CLK=>nx34513);
   reg_label_10_input_state_machine_9 : dffr port map ( Q=>
      label_10_input_state_machine_9, QB=>OPEN, D=>nx18883, CLK=>clk, R=>rst
   );
   ix8417 : xnor2 port map ( Y=>nx8416, A0=>nx8406, A1=>nx27724);
   ix8407 : oai22 port map ( Y=>nx8406, A0=>nx27619, A1=>nx27713, B0=>
      nx27723, B1=>nx27560);
   ix27620 : aoi22 port map ( Y=>nx27619, A0=>label_10_output(7), A1=>
      booth_booth_integration_output_9_7, B0=>nx8342, B1=>nx13187);
   labelsregfile_label10_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_10_output(7), QB=>OPEN, D=>nx18853, CLK=>clk, R=>rst);
   lat_label_10_input_7 : latch port map ( Q=>label_10_input_7, D=>nx8356, 
      CLK=>nx34513);
   reg_label_10_input_state_machine_7 : dffr port map ( Q=>
      label_10_input_state_machine_7, QB=>OPEN, D=>nx18843, CLK=>clk, R=>rst
   );
   ix8353 : xnor2 port map ( Y=>nx8352, A0=>nx8342, A1=>nx27709);
   ix8343 : oai22 port map ( Y=>nx8342, A0=>nx27630, A1=>nx27698, B0=>
      nx27708, B1=>nx27562);
   ix27631 : aoi22 port map ( Y=>nx27630, A0=>label_10_output(5), A1=>
      booth_booth_integration_output_9_5, B0=>nx8278, B1=>nx13183);
   labelsregfile_label10_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_10_output(5), QB=>OPEN, D=>nx18813, CLK=>clk, R=>rst);
   lat_label_10_input_5 : latch port map ( Q=>label_10_input_5, D=>nx8292, 
      CLK=>nx34513);
   reg_label_10_input_state_machine_5 : dffr port map ( Q=>
      label_10_input_state_machine_5, QB=>OPEN, D=>nx18803, CLK=>clk, R=>rst
   );
   ix8289 : xnor2 port map ( Y=>nx8288, A0=>nx8278, A1=>nx27694);
   ix8279 : oai22 port map ( Y=>nx8278, A0=>nx27641, A1=>nx27683, B0=>
      nx27693, B1=>nx27564);
   ix27642 : aoi22 port map ( Y=>nx27641, A0=>label_10_output(3), A1=>
      booth_booth_integration_output_9_3, B0=>nx8214, B1=>nx13179);
   labelsregfile_label10_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_10_output(3), QB=>OPEN, D=>nx18773, CLK=>clk, R=>rst);
   lat_label_10_input_3 : latch port map ( Q=>label_10_input_3, D=>nx8228, 
      CLK=>nx34511);
   reg_label_10_input_state_machine_3 : dffr port map ( Q=>
      label_10_input_state_machine_3, QB=>OPEN, D=>nx18763, CLK=>clk, R=>rst
   );
   ix8225 : xnor2 port map ( Y=>nx8224, A0=>nx8214, A1=>nx27679);
   ix8215 : oai22 port map ( Y=>nx8214, A0=>nx27652, A1=>nx27668, B0=>
      nx27678, B1=>nx27566);
   ix27653 : aoi32 port map ( Y=>nx27652, A0=>label_10_output(0), A1=>
      nx35759, A2=>nx13175, B0=>label_10_output(1), B1=>
      booth_booth_integration_output_9_1);
   labelsregfile_label10_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_10_output(1), QB=>OPEN, D=>nx18733, CLK=>clk, R=>rst);
   lat_label_10_input_1 : latch port map ( Q=>label_10_input_1, D=>nx8164, 
      CLK=>nx34511);
   reg_label_10_input_state_machine_1 : dffr port map ( Q=>
      label_10_input_state_machine_1, QB=>OPEN, D=>nx18723, CLK=>clk, R=>rst
   );
   ix8161 : xor2 port map ( Y=>nx8160, A0=>nx27663, A1=>nx27665);
   ix27664 : nand02 port map ( Y=>nx27663, A0=>label_10_output(0), A1=>
      nx35759);
   ix27666 : xnor2 port map ( Y=>nx27665, A0=>
      booth_booth_integration_output_9_1, A1=>label_10_output(1));
   labelsregfile_label10_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_10_output(2), QB=>nx27678, D=>nx18753, CLK=>clk, R=>rst);
   lat_label_10_input_2 : latch port map ( Q=>label_10_input_2, D=>nx8196, 
      CLK=>nx34511);
   reg_label_10_input_state_machine_2 : dffr port map ( Q=>
      label_10_input_state_machine_2, QB=>OPEN, D=>nx18743, CLK=>clk, R=>rst
   );
   ix8193 : xor2 port map ( Y=>nx8192, A0=>nx27652, A1=>nx27668);
   ix27680 : xnor2 port map ( Y=>nx27679, A0=>
      booth_booth_integration_output_9_3, A1=>label_10_output(3));
   labelsregfile_label10_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_10_output(4), QB=>nx27693, D=>nx18793, CLK=>clk, R=>rst);
   lat_label_10_input_4 : latch port map ( Q=>label_10_input_4, D=>nx8260, 
      CLK=>nx34511);
   reg_label_10_input_state_machine_4 : dffr port map ( Q=>
      label_10_input_state_machine_4, QB=>OPEN, D=>nx18783, CLK=>clk, R=>rst
   );
   ix8257 : xor2 port map ( Y=>nx8256, A0=>nx27641, A1=>nx27683);
   ix27695 : xnor2 port map ( Y=>nx27694, A0=>
      booth_booth_integration_output_9_5, A1=>label_10_output(5));
   labelsregfile_label10_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_10_output(6), QB=>nx27708, D=>nx18833, CLK=>clk, R=>rst);
   lat_label_10_input_6 : latch port map ( Q=>label_10_input_6, D=>nx8324, 
      CLK=>nx34513);
   reg_label_10_input_state_machine_6 : dffr port map ( Q=>
      label_10_input_state_machine_6, QB=>OPEN, D=>nx18823, CLK=>clk, R=>rst
   );
   ix8321 : xor2 port map ( Y=>nx8320, A0=>nx27630, A1=>nx27698);
   ix27710 : xnor2 port map ( Y=>nx27709, A0=>
      booth_booth_integration_output_9_7, A1=>label_10_output(7));
   labelsregfile_label10_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_10_output(8), QB=>nx27723, D=>nx18873, CLK=>clk, R=>rst);
   lat_label_10_input_8 : latch port map ( Q=>label_10_input_8, D=>nx8388, 
      CLK=>nx34513);
   reg_label_10_input_state_machine_8 : dffr port map ( Q=>
      label_10_input_state_machine_8, QB=>OPEN, D=>nx18863, CLK=>clk, R=>rst
   );
   ix8385 : xor2 port map ( Y=>nx8384, A0=>nx27619, A1=>nx27713);
   ix27725 : xnor2 port map ( Y=>nx27724, A0=>
      booth_booth_integration_output_9_9, A1=>label_10_output(9));
   labelsregfile_label10_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_10_output(10), QB=>nx27738, D=>nx18913, CLK=>clk, R=>rst);
   lat_label_10_input_10 : latch port map ( Q=>label_10_input_10, D=>nx8452, 
      CLK=>nx34513);
   reg_label_10_input_state_machine_10 : dffr port map ( Q=>
      label_10_input_state_machine_10, QB=>OPEN, D=>nx18903, CLK=>clk, R=>
      rst);
   ix8449 : xor2 port map ( Y=>nx8448, A0=>nx27608, A1=>nx27728);
   ix27740 : xnor2 port map ( Y=>nx27739, A0=>
      booth_booth_integration_output_9_11, A1=>label_10_output(11));
   labelsregfile_label10_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_10_output(12), QB=>nx27753, D=>nx18953, CLK=>clk, R=>rst);
   lat_label_10_input_12 : latch port map ( Q=>label_10_input_12, D=>nx8516, 
      CLK=>nx34515);
   reg_label_10_input_state_machine_12 : dffr port map ( Q=>
      label_10_input_state_machine_12, QB=>OPEN, D=>nx18943, CLK=>clk, R=>
      rst);
   ix8513 : xor2 port map ( Y=>nx8512, A0=>nx27597, A1=>nx27743);
   ix27755 : xnor2 port map ( Y=>nx27754, A0=>
      booth_booth_integration_output_9_13, A1=>label_10_output(13));
   ix19284 : oai21 port map ( Y=>nx19283, A0=>nx27763, A1=>nx34747, B0=>
      nx27765);
   max_calc_reg_comparator_fifth_inp1_14 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_14, QB=>nx27763, D=>nx19283, CLK=>clk);
   labelsregfile_label9_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_9_output(14), QB=>nx27949, D=>nx19273, CLK=>clk, R=>rst);
   lat_label_9_input_14 : latch port map ( Q=>label_9_input_14, D=>nx9024, 
      CLK=>nx34519);
   reg_label_9_input_state_machine_14 : dffr port map ( Q=>
      label_9_input_state_machine_14, QB=>OPEN, D=>nx19003, CLK=>clk, R=>rst
   );
   ix9021 : xor2 port map ( Y=>nx9020, A0=>nx27775, A1=>nx27947);
   ix27776 : aoi22 port map ( Y=>nx27775, A0=>label_9_output(13), A1=>
      booth_booth_integration_output_8_13, B0=>nx8984, B1=>nx13215);
   labelsregfile_label9_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_9_output(13), QB=>OPEN, D=>nx19263, CLK=>clk, R=>rst);
   lat_label_9_input_13 : latch port map ( Q=>label_9_input_13, D=>nx8998, 
      CLK=>nx34519);
   reg_label_9_input_state_machine_13 : dffr port map ( Q=>
      label_9_input_state_machine_13, QB=>OPEN, D=>nx19253, CLK=>clk, R=>rst
   );
   ix8995 : xnor2 port map ( Y=>nx8994, A0=>nx8984, A1=>nx27943);
   ix8985 : oai22 port map ( Y=>nx8984, A0=>nx27786, A1=>nx27932, B0=>
      nx27942, B1=>nx27117);
   ix27787 : aoi22 port map ( Y=>nx27786, A0=>label_9_output(11), A1=>
      booth_booth_integration_output_8_11, B0=>nx8920, B1=>nx13213);
   labelsregfile_label9_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_9_output(11), QB=>OPEN, D=>nx19223, CLK=>clk, R=>rst);
   lat_label_9_input_11 : latch port map ( Q=>label_9_input_11, D=>nx8934, 
      CLK=>nx34517);
   reg_label_9_input_state_machine_11 : dffr port map ( Q=>
      label_9_input_state_machine_11, QB=>OPEN, D=>nx19213, CLK=>clk, R=>rst
   );
   ix8931 : xnor2 port map ( Y=>nx8930, A0=>nx8920, A1=>nx27928);
   ix8921 : oai22 port map ( Y=>nx8920, A0=>nx27797, A1=>nx27917, B0=>
      nx27927, B1=>nx27119);
   ix27798 : aoi22 port map ( Y=>nx27797, A0=>label_9_output(9), A1=>
      booth_booth_integration_output_8_9, B0=>nx8856, B1=>nx13211);
   labelsregfile_label9_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_9_output(9), QB=>OPEN, D=>nx19183, CLK=>clk, R=>rst);
   lat_label_9_input_9 : latch port map ( Q=>label_9_input_9, D=>nx8870, CLK
      =>nx34517);
   reg_label_9_input_state_machine_9 : dffr port map ( Q=>
      label_9_input_state_machine_9, QB=>OPEN, D=>nx19173, CLK=>clk, R=>rst
   );
   ix8867 : xnor2 port map ( Y=>nx8866, A0=>nx8856, A1=>nx27913);
   ix8857 : oai22 port map ( Y=>nx8856, A0=>nx27808, A1=>nx27902, B0=>
      nx27912, B1=>nx27121);
   ix27809 : aoi22 port map ( Y=>nx27808, A0=>label_9_output(7), A1=>
      booth_booth_integration_output_8_7, B0=>nx8792, B1=>nx13207);
   labelsregfile_label9_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_9_output(7), QB=>OPEN, D=>nx19143, CLK=>clk, R=>rst);
   lat_label_9_input_7 : latch port map ( Q=>label_9_input_7, D=>nx8806, CLK
      =>nx34517);
   reg_label_9_input_state_machine_7 : dffr port map ( Q=>
      label_9_input_state_machine_7, QB=>OPEN, D=>nx19133, CLK=>clk, R=>rst
   );
   ix8803 : xnor2 port map ( Y=>nx8802, A0=>nx8792, A1=>nx27898);
   ix8793 : oai22 port map ( Y=>nx8792, A0=>nx27819, A1=>nx27887, B0=>
      nx27897, B1=>nx27123);
   ix27820 : aoi22 port map ( Y=>nx27819, A0=>label_9_output(5), A1=>
      booth_booth_integration_output_8_5, B0=>nx8728, B1=>nx13204);
   labelsregfile_label9_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_9_output(5), QB=>OPEN, D=>nx19103, CLK=>clk, R=>rst);
   lat_label_9_input_5 : latch port map ( Q=>label_9_input_5, D=>nx8742, CLK
      =>nx34517);
   reg_label_9_input_state_machine_5 : dffr port map ( Q=>
      label_9_input_state_machine_5, QB=>OPEN, D=>nx19093, CLK=>clk, R=>rst
   );
   ix8739 : xnor2 port map ( Y=>nx8738, A0=>nx8728, A1=>nx27883);
   ix8729 : oai22 port map ( Y=>nx8728, A0=>nx27830, A1=>nx27872, B0=>
      nx27882, B1=>nx27125);
   ix27831 : aoi22 port map ( Y=>nx27830, A0=>label_9_output(3), A1=>
      booth_booth_integration_output_8_3, B0=>nx8664, B1=>nx13202);
   labelsregfile_label9_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_9_output(3), QB=>OPEN, D=>nx19063, CLK=>clk, R=>rst);
   lat_label_9_input_3 : latch port map ( Q=>label_9_input_3, D=>nx8678, CLK
      =>nx34515);
   reg_label_9_input_state_machine_3 : dffr port map ( Q=>
      label_9_input_state_machine_3, QB=>OPEN, D=>nx19053, CLK=>clk, R=>rst
   );
   ix8675 : xnor2 port map ( Y=>nx8674, A0=>nx8664, A1=>nx27868);
   ix8665 : oai22 port map ( Y=>nx8664, A0=>nx27841, A1=>nx27857, B0=>
      nx27867, B1=>nx27127);
   ix27842 : aoi32 port map ( Y=>nx27841, A0=>label_9_output(0), A1=>nx35755, 
      A2=>nx13200, B0=>label_9_output(1), B1=>
      booth_booth_integration_output_8_1);
   labelsregfile_label9_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_9_output(1), QB=>OPEN, D=>nx19023, CLK=>clk, R=>rst);
   lat_label_9_input_1 : latch port map ( Q=>label_9_input_1, D=>nx8614, CLK
      =>nx34515);
   reg_label_9_input_state_machine_1 : dffr port map ( Q=>
      label_9_input_state_machine_1, QB=>OPEN, D=>nx19013, CLK=>clk, R=>rst
   );
   ix8611 : xor2 port map ( Y=>nx8610, A0=>nx27852, A1=>nx27854);
   ix27853 : nand02 port map ( Y=>nx27852, A0=>label_9_output(0), A1=>
      nx35755);
   ix27855 : xnor2 port map ( Y=>nx27854, A0=>
      booth_booth_integration_output_8_1, A1=>label_9_output(1));
   labelsregfile_label9_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_9_output(2), QB=>nx27867, D=>nx19043, CLK=>clk, R=>rst);
   lat_label_9_input_2 : latch port map ( Q=>label_9_input_2, D=>nx8646, CLK
      =>nx34515);
   reg_label_9_input_state_machine_2 : dffr port map ( Q=>
      label_9_input_state_machine_2, QB=>OPEN, D=>nx19033, CLK=>clk, R=>rst
   );
   ix8643 : xor2 port map ( Y=>nx8642, A0=>nx27841, A1=>nx27857);
   ix27869 : xnor2 port map ( Y=>nx27868, A0=>
      booth_booth_integration_output_8_3, A1=>label_9_output(3));
   labelsregfile_label9_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_9_output(4), QB=>nx27882, D=>nx19083, CLK=>clk, R=>rst);
   lat_label_9_input_4 : latch port map ( Q=>label_9_input_4, D=>nx8710, CLK
      =>nx34515);
   reg_label_9_input_state_machine_4 : dffr port map ( Q=>
      label_9_input_state_machine_4, QB=>OPEN, D=>nx19073, CLK=>clk, R=>rst
   );
   ix8707 : xor2 port map ( Y=>nx8706, A0=>nx27830, A1=>nx27872);
   ix27884 : xnor2 port map ( Y=>nx27883, A0=>
      booth_booth_integration_output_8_5, A1=>label_9_output(5));
   labelsregfile_label9_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_9_output(6), QB=>nx27897, D=>nx19123, CLK=>clk, R=>rst);
   lat_label_9_input_6 : latch port map ( Q=>label_9_input_6, D=>nx8774, CLK
      =>nx34517);
   reg_label_9_input_state_machine_6 : dffr port map ( Q=>
      label_9_input_state_machine_6, QB=>OPEN, D=>nx19113, CLK=>clk, R=>rst
   );
   ix8771 : xor2 port map ( Y=>nx8770, A0=>nx27819, A1=>nx27887);
   ix27899 : xnor2 port map ( Y=>nx27898, A0=>
      booth_booth_integration_output_8_7, A1=>label_9_output(7));
   labelsregfile_label9_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_9_output(8), QB=>nx27912, D=>nx19163, CLK=>clk, R=>rst);
   lat_label_9_input_8 : latch port map ( Q=>label_9_input_8, D=>nx8838, CLK
      =>nx34517);
   reg_label_9_input_state_machine_8 : dffr port map ( Q=>
      label_9_input_state_machine_8, QB=>OPEN, D=>nx19153, CLK=>clk, R=>rst
   );
   ix8835 : xor2 port map ( Y=>nx8834, A0=>nx27808, A1=>nx27902);
   ix27914 : xnor2 port map ( Y=>nx27913, A0=>
      booth_booth_integration_output_8_9, A1=>label_9_output(9));
   labelsregfile_label9_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_9_output(10), QB=>nx27927, D=>nx19203, CLK=>clk, R=>rst);
   lat_label_9_input_10 : latch port map ( Q=>label_9_input_10, D=>nx8902, 
      CLK=>nx34517);
   reg_label_9_input_state_machine_10 : dffr port map ( Q=>
      label_9_input_state_machine_10, QB=>OPEN, D=>nx19193, CLK=>clk, R=>rst
   );
   ix8899 : xor2 port map ( Y=>nx8898, A0=>nx27797, A1=>nx27917);
   ix27929 : xnor2 port map ( Y=>nx27928, A0=>
      booth_booth_integration_output_8_11, A1=>label_9_output(11));
   labelsregfile_label9_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_9_output(12), QB=>nx27942, D=>nx19243, CLK=>clk, R=>rst);
   lat_label_9_input_12 : latch port map ( Q=>label_9_input_12, D=>nx8966, 
      CLK=>nx34519);
   reg_label_9_input_state_machine_12 : dffr port map ( Q=>
      label_9_input_state_machine_12, QB=>OPEN, D=>nx19233, CLK=>clk, R=>rst
   );
   ix8963 : xor2 port map ( Y=>nx8962, A0=>nx27786, A1=>nx27932);
   ix27944 : xnor2 port map ( Y=>nx27943, A0=>
      booth_booth_integration_output_8_13, A1=>label_9_output(13));
   ix9399 : oai22 port map ( Y=>nx9398, A0=>nx27952, A1=>nx27965, B0=>
      max_calc_comparator_fifth_inp2_13, B1=>nx27960);
   ix19294 : oai21 port map ( Y=>nx19293, A0=>nx27956, A1=>nx34749, B0=>
      nx27958);
   max_calc_reg_comparator_fifth_inp2_13 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_13, QB=>nx27956, D=>nx19293, CLK=>clk);
   ix27959 : nand03 port map ( Y=>nx27958, A0=>label_10_output(13), A1=>
      nx34737, A2=>nx34749);
   max_calc_reg_comparator_fifth_inp1_13 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_13, QB=>nx27960, D=>nx19303, CLK=>clk);
   ix19304 : oai21 port map ( Y=>nx19303, A0=>nx27960, A1=>nx34749, B0=>
      nx27963);
   ix27964 : nand03 port map ( Y=>nx27963, A0=>label_9_output(13), A1=>
      nx34739, A2=>nx34749);
   ix27966 : aoi22 port map ( Y=>nx27965, A0=>nx27967, A1=>
      max_calc_comparator_fifth_inp1_12, B0=>nx9080, B1=>nx9382);
   max_calc_reg_comparator_fifth_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx27967, D=>nx19313, CLK=>clk);
   ix19314 : oai21 port map ( Y=>nx19313, A0=>nx27967, A1=>nx34749, B0=>
      nx27970);
   ix19324 : oai21 port map ( Y=>nx19323, A0=>nx27974, A1=>nx34751, B0=>
      nx27976);
   max_calc_reg_comparator_fifth_inp1_12 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_12, QB=>nx27974, D=>nx19323, CLK=>clk);
   ix9383 : oai22 port map ( Y=>nx9382, A0=>nx27980, A1=>nx27993, B0=>
      max_calc_comparator_fifth_inp2_11, B1=>nx27988);
   ix19334 : oai21 port map ( Y=>nx19333, A0=>nx27984, A1=>nx34751, B0=>
      nx27986);
   max_calc_reg_comparator_fifth_inp2_11 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_11, QB=>nx27984, D=>nx19333, CLK=>clk);
   ix27987 : nand03 port map ( Y=>nx27986, A0=>label_10_output(11), A1=>
      nx34739, A2=>nx34751);
   max_calc_reg_comparator_fifth_inp1_11 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_11, QB=>nx27988, D=>nx19343, CLK=>clk);
   ix19344 : oai21 port map ( Y=>nx19343, A0=>nx27988, A1=>nx34751, B0=>
      nx27991);
   ix27992 : nand03 port map ( Y=>nx27991, A0=>label_9_output(11), A1=>
      nx34739, A2=>nx34751);
   ix27994 : aoi22 port map ( Y=>nx27993, A0=>nx27995, A1=>
      max_calc_comparator_fifth_inp1_10, B0=>nx9116, B1=>nx9366);
   max_calc_reg_comparator_fifth_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx27995, D=>nx19353, CLK=>clk);
   ix19354 : oai21 port map ( Y=>nx19353, A0=>nx27995, A1=>nx34751, B0=>
      nx27998);
   ix19364 : oai21 port map ( Y=>nx19363, A0=>nx28002, A1=>nx34753, B0=>
      nx28004);
   max_calc_reg_comparator_fifth_inp1_10 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_10, QB=>nx28002, D=>nx19363, CLK=>clk);
   ix9367 : oai22 port map ( Y=>nx9366, A0=>nx28008, A1=>nx28021, B0=>
      max_calc_comparator_fifth_inp2_9, B1=>nx28016);
   ix19374 : oai21 port map ( Y=>nx19373, A0=>nx28012, A1=>nx34753, B0=>
      nx28014);
   max_calc_reg_comparator_fifth_inp2_9 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_9, QB=>nx28012, D=>nx19373, CLK=>clk);
   ix28015 : nand03 port map ( Y=>nx28014, A0=>label_10_output(9), A1=>
      nx34741, A2=>nx34753);
   max_calc_reg_comparator_fifth_inp1_9 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_9, QB=>nx28016, D=>nx19383, CLK=>clk);
   ix19384 : oai21 port map ( Y=>nx19383, A0=>nx28016, A1=>nx34753, B0=>
      nx28019);
   ix28020 : nand03 port map ( Y=>nx28019, A0=>label_9_output(9), A1=>
      nx34741, A2=>nx34753);
   ix28022 : aoi22 port map ( Y=>nx28021, A0=>nx28023, A1=>
      max_calc_comparator_fifth_inp1_8, B0=>nx9152, B1=>nx9350);
   max_calc_reg_comparator_fifth_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx28023, D=>nx19393, CLK=>clk);
   ix19394 : oai21 port map ( Y=>nx19393, A0=>nx28023, A1=>nx34755, B0=>
      nx28026);
   ix19404 : oai21 port map ( Y=>nx19403, A0=>nx28030, A1=>nx34755, B0=>
      nx28032);
   max_calc_reg_comparator_fifth_inp1_8 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_8, QB=>nx28030, D=>nx19403, CLK=>clk);
   ix9351 : oai22 port map ( Y=>nx9350, A0=>nx28036, A1=>nx28049, B0=>
      max_calc_comparator_fifth_inp2_7, B1=>nx28044);
   ix19414 : oai21 port map ( Y=>nx19413, A0=>nx28040, A1=>nx34755, B0=>
      nx28042);
   max_calc_reg_comparator_fifth_inp2_7 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_7, QB=>nx28040, D=>nx19413, CLK=>clk);
   ix28043 : nand03 port map ( Y=>nx28042, A0=>label_10_output(7), A1=>
      nx34741, A2=>nx34755);
   max_calc_reg_comparator_fifth_inp1_7 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_7, QB=>nx28044, D=>nx19423, CLK=>clk);
   ix19424 : oai21 port map ( Y=>nx19423, A0=>nx28044, A1=>nx34755, B0=>
      nx28047);
   ix28048 : nand03 port map ( Y=>nx28047, A0=>label_9_output(7), A1=>
      nx34741, A2=>nx34757);
   ix28050 : aoi22 port map ( Y=>nx28049, A0=>nx28051, A1=>
      max_calc_comparator_fifth_inp1_6, B0=>nx9188, B1=>nx9334);
   max_calc_reg_comparator_fifth_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx28051, D=>nx19433, CLK=>clk);
   ix19434 : oai21 port map ( Y=>nx19433, A0=>nx28051, A1=>nx34757, B0=>
      nx28054);
   ix19444 : oai21 port map ( Y=>nx19443, A0=>nx28058, A1=>nx34757, B0=>
      nx28060);
   max_calc_reg_comparator_fifth_inp1_6 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_6, QB=>nx28058, D=>nx19443, CLK=>clk);
   ix9335 : oai22 port map ( Y=>nx9334, A0=>nx28064, A1=>nx28077, B0=>
      max_calc_comparator_fifth_inp2_5, B1=>nx28072);
   ix19454 : oai21 port map ( Y=>nx19453, A0=>nx28068, A1=>nx34757, B0=>
      nx28070);
   max_calc_reg_comparator_fifth_inp2_5 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_5, QB=>nx28068, D=>nx19453, CLK=>clk);
   ix28071 : nand03 port map ( Y=>nx28070, A0=>label_10_output(5), A1=>
      nx34743, A2=>nx34757);
   max_calc_reg_comparator_fifth_inp1_5 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_5, QB=>nx28072, D=>nx19463, CLK=>clk);
   ix19464 : oai21 port map ( Y=>nx19463, A0=>nx28072, A1=>nx34759, B0=>
      nx28075);
   ix28076 : nand03 port map ( Y=>nx28075, A0=>label_9_output(5), A1=>
      nx34743, A2=>nx34759);
   ix28078 : aoi22 port map ( Y=>nx28077, A0=>nx28079, A1=>
      max_calc_comparator_fifth_inp1_4, B0=>nx9224, B1=>nx9318);
   max_calc_reg_comparator_fifth_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx28079, D=>nx19473, CLK=>clk);
   ix19474 : oai21 port map ( Y=>nx19473, A0=>nx28079, A1=>nx34759, B0=>
      nx28082);
   ix19484 : oai21 port map ( Y=>nx19483, A0=>nx28086, A1=>nx34759, B0=>
      nx28088);
   max_calc_reg_comparator_fifth_inp1_4 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_4, QB=>nx28086, D=>nx19483, CLK=>clk);
   ix9319 : oai22 port map ( Y=>nx9318, A0=>nx28092, A1=>nx28105, B0=>
      max_calc_comparator_fifth_inp2_3, B1=>nx28100);
   ix19494 : oai21 port map ( Y=>nx19493, A0=>nx28096, A1=>nx34759, B0=>
      nx28098);
   max_calc_reg_comparator_fifth_inp2_3 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_3, QB=>nx28096, D=>nx19493, CLK=>clk);
   ix28099 : nand03 port map ( Y=>nx28098, A0=>label_10_output(3), A1=>
      nx34743, A2=>nx34761);
   max_calc_reg_comparator_fifth_inp1_3 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_3, QB=>nx28100, D=>nx19503, CLK=>clk);
   ix19504 : oai21 port map ( Y=>nx19503, A0=>nx28100, A1=>nx34761, B0=>
      nx28103);
   ix28104 : nand03 port map ( Y=>nx28103, A0=>label_9_output(3), A1=>
      nx34743, A2=>nx34761);
   ix28106 : aoi22 port map ( Y=>nx28105, A0=>nx28107, A1=>
      max_calc_comparator_fifth_inp1_2, B0=>nx9260, B1=>nx9302);
   max_calc_reg_comparator_fifth_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx28107, D=>nx19513, CLK=>clk);
   ix19514 : oai21 port map ( Y=>nx19513, A0=>nx28107, A1=>nx34761, B0=>
      nx28110);
   ix19524 : oai21 port map ( Y=>nx19523, A0=>nx28114, A1=>nx34761, B0=>
      nx28116);
   max_calc_reg_comparator_fifth_inp1_2 : dff port map ( Q=>
      max_calc_comparator_fifth_inp1_2, QB=>nx28114, D=>nx19523, CLK=>clk);
   ix9303 : oai21 port map ( Y=>nx9302, A0=>max_calc_comparator_fifth_inp2_1, 
      A1=>nx28126, B0=>nx28131);
   ix19534 : oai21 port map ( Y=>nx19533, A0=>nx28122, A1=>nx34763, B0=>
      nx28124);
   max_calc_reg_comparator_fifth_inp2_1 : dff port map ( Q=>
      max_calc_comparator_fifth_inp2_1, QB=>nx28122, D=>nx19533, CLK=>clk);
   ix28125 : nand03 port map ( Y=>nx28124, A0=>label_10_output(1), A1=>
      nx34745, A2=>nx34763);
   max_calc_reg_comparator_fifth_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx28126, D=>nx19543, CLK=>clk);
   ix19544 : oai21 port map ( Y=>nx19543, A0=>nx28126, A1=>nx34763, B0=>
      nx28129);
   ix28130 : nand03 port map ( Y=>nx28129, A0=>label_9_output(1), A1=>
      nx34745, A2=>nx34763);
   ix28132 : oai21 port map ( Y=>nx28131, A0=>nx27133, A1=>
      max_calc_comparator_fifth_inp1_0, B0=>nx9278);
   ix19584 : oai21 port map ( Y=>nx19583, A0=>nx28137, A1=>nx34763, B0=>
      nx28139);
   max_calc_reg_comparator_fifth_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx28137, D=>nx19583, CLK=>clk);
   ix28140 : nand03 port map ( Y=>nx28139, A0=>label_10_output(15), A1=>
      nx34745, A2=>nx34763);
   labelsregfile_label10_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_10_output(15), QB=>OPEN, D=>nx19573, CLK=>clk, R=>rst);
   lat_label_10_input_15 : latch port map ( Q=>label_10_input_15, D=>nx9428, 
      CLK=>nx34519);
   reg_label_10_input_state_machine_15 : dffr port map ( Q=>
      label_10_input_state_machine_15, QB=>OPEN, D=>nx19563, CLK=>clk, R=>
      rst);
   ix9425 : xnor2 port map ( Y=>nx9424, A0=>nx9420, A1=>nx28150);
   ix9421 : oai22 port map ( Y=>nx9420, A0=>nx27586, A1=>nx27758, B0=>
      nx27760, B1=>nx27554);
   ix19614 : oai21 port map ( Y=>nx19613, A0=>nx28155, A1=>nx34763, B0=>
      nx28157);
   max_calc_reg_comparator_fifth_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx28155, D=>nx19613, CLK=>clk);
   ix28158 : nand03 port map ( Y=>nx28157, A0=>label_9_output(15), A1=>
      nx34745, A2=>nx34765);
   labelsregfile_label9_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_9_output(15), QB=>OPEN, D=>nx19603, CLK=>clk, R=>rst);
   lat_label_9_input_15 : latch port map ( Q=>label_9_input_15, D=>nx9468, 
      CLK=>nx34519);
   reg_label_9_input_state_machine_15 : dffr port map ( Q=>
      label_9_input_state_machine_15, QB=>OPEN, D=>nx19593, CLK=>clk, R=>rst
   );
   ix9465 : xnor2 port map ( Y=>nx9464, A0=>nx9460, A1=>nx28168);
   ix9461 : oai22 port map ( Y=>nx9460, A0=>nx27775, A1=>nx27947, B0=>
      nx27949, B1=>nx27115);
   max_calc_reg_comparator_first_inp2_0 : dff port map ( Q=>
      max_calc_comparator_first_inp2_0, QB=>nx33288, D=>nx25473, CLK=>clk);
   labelsregfile_label2_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_2_output(0), QB=>OPEN, D=>nx16373, CLK=>clk, R=>rst);
   lat_label_2_input_0 : latch port map ( Q=>label_2_input_0, D=>nx4420, CLK
      =>nx34519);
   ix4421 : oai21 port map ( Y=>nx4420, A0=>nx28183, A1=>nx34419, B0=>
      nx28187);
   reg_label_2_input_state_machine_0 : dffr port map ( Q=>
      label_2_input_state_machine_0, QB=>nx28183, D=>nx16363, CLK=>clk, R=>
      rst);
   ix28188 : oai21 port map ( Y=>nx28187, A0=>nx35727, A1=>label_2_output(0), 
      B0=>nx4408);
   booth_booth_integrtaion_1_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_1, QB=>OPEN, D=>nx16343, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_2, QB=>nx28608, D=>nx16333, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_3, QB=>OPEN, D=>nx16323, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_4, QB=>nx28606, D=>nx16313, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_5, QB=>OPEN, D=>nx16303, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_6, QB=>nx28604, D=>nx16293, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_7, QB=>OPEN, D=>nx16283, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_8, QB=>nx28602, D=>nx16273, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_9, QB=>OPEN, D=>nx16263, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_10, QB=>nx28600, D=>nx16253, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_11, QB=>OPEN, D=>nx16243, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_12, QB=>nx28598, D=>nx16233, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_13, QB=>OPEN, D=>nx16223, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_14, QB=>nx28596, D=>nx16213, CLK=>clk, 
      R=>rst);
   ix28237 : aoi22 port map ( Y=>nx28236, A0=>mdr_data_out(15), A1=>nx34635, 
      B0=>nx4206, B1=>nx4212);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_reg_output_0, QB=>OPEN, 
      D=>nx15853, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_0, QB=>OPEN, D=>nx15839, CLK
      =>clk, S=>nx34475);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_reg_output_9, QB=>OPEN, 
      D=>nx16033, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_9, QB=>OPEN, D=>nx16023, CLK
      =>clk, R=>nx34473);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_8, QB=>OPEN, 
      D=>nx16013, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_8, QB=>OPEN, D=>nx16003, CLK
      =>clk, R=>nx34473);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_7, QB=>OPEN, 
      D=>nx15993, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_7, QB=>OPEN, D=>nx15983, CLK
      =>clk, R=>nx34473);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_6, QB=>OPEN, 
      D=>nx15973, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_6, QB=>OPEN, D=>nx15963, CLK
      =>clk, R=>nx34473);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_5, QB=>OPEN, 
      D=>nx15953, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_5, QB=>OPEN, D=>nx15943, CLK
      =>clk, R=>nx34473);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_4, QB=>OPEN, 
      D=>nx15933, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_4, QB=>OPEN, D=>nx15923, CLK
      =>clk, R=>nx34473);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_3, QB=>OPEN, 
      D=>nx15913, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_3, QB=>OPEN, D=>nx15903, CLK
      =>clk, R=>nx34473);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_2, QB=>OPEN, 
      D=>nx15893, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_2, QB=>OPEN, D=>nx15883, CLK
      =>clk, R=>nx34471);
   booth_booth_integrtaion_1_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_1_shift_Reg_output_1, QB=>OPEN, 
      D=>nx15873, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_1_shift_Reg_count_1, QB=>OPEN, D=>nx15863, CLK
      =>clk, R=>nx34471);
   ix15834 : nand02 port map ( Y=>nx15833, A0=>nx35815, A1=>nx34621);
   booth_booth_integrtaion_1_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx28283, D=>nx15833, CLK=>clk, S=>nx34471);
   ix4207 : nand02 port map ( Y=>nx4206, A0=>nx28304, A1=>nx28316);
   ix28305 : oai21 port map ( Y=>nx28304, A0=>nx34649, A1=>nx34643, B0=>
      mdr_data_out(32));
   ix16044 : oai21 port map ( Y=>nx16043, A0=>nx28309, A1=>nx35373, B0=>
      nx28311);
   booth_booth_integrtaion_1_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx28309, D=>nx16043, CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx28313, D=>nx16353, CLK=>clk, R=>rst);
   ix28321 : xnor2 port map ( Y=>nx28320, A0=>nx3676, A1=>nx13017);
   ix16184 : oai21 port map ( Y=>nx16183, A0=>nx28326, A1=>nx35373, B0=>
      nx28328);
   booth_booth_integrtaion_1_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_17, QB=>nx28326, D=>nx16183, 
      CLK=>clk, R=>rst);
   ix28329 : nand03 port map ( Y=>nx28328, A0=>nx35381, A1=>nx4184, A2=>
      nx36077);
   ix4185 : xnor2 port map ( Y=>nx4184, A0=>nx28331, A1=>nx13018);
   ix28332 : aoi22 port map ( Y=>nx28331, A0=>
      booth_booth_integrtaion_1_booth_output_17, A1=>nx3700, B0=>nx3676, B1
      =>nx13017);
   ix3685 : nand02 port map ( Y=>nx3684, A0=>mdr_data_out(33), A1=>
      mdr_data_out(32));
   ix28336 : or02 port map ( Y=>nx28335, A0=>mdr_data_out(32), A1=>
      mdr_data_out(33));
   ix28342 : xnor2 port map ( Y=>nx28341, A0=>nx3728, A1=>nx13019);
   ix3729 : oai22 port map ( Y=>nx3728, A0=>nx28331, A1=>nx28344, B0=>
      nx28351, B1=>nx35385);
   ix28347 : aoi32 port map ( Y=>nx28346, A0=>nx3710, A1=>nx34649, A2=>
      nx28349, B0=>mdr_data_out(34), B1=>nx34643);
   ix3711 : oai21 port map ( Y=>nx3710, A0=>mdr_data_out(32), A1=>
      mdr_data_out(33), B0=>mdr_data_out(34));
   booth_booth_integrtaion_1_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_18, QB=>nx28351, D=>nx16173, 
      CLK=>clk, R=>rst);
   ix16164 : oai21 port map ( Y=>nx16163, A0=>nx28356, A1=>nx35373, B0=>
      nx28358);
   booth_booth_integrtaion_1_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_19, QB=>nx28356, D=>nx16163, 
      CLK=>clk, R=>rst);
   ix28359 : nand03 port map ( Y=>nx28358, A0=>nx35381, A1=>nx4160, A2=>
      nx36077);
   ix4161 : xnor2 port map ( Y=>nx4160, A0=>nx28361, A1=>nx13021);
   ix28362 : aoi22 port map ( Y=>nx28361, A0=>
      booth_booth_integrtaion_1_booth_output_19, A1=>nx3748, B0=>nx3728, B1
      =>nx13019);
   ix28365 : nor02ii port map ( Y=>nx28364, A0=>nx3714, A1=>mdr_data_out(35)
   );
   ix3715 : nor03_2x port map ( Y=>nx3714, A0=>mdr_data_out(34), A1=>
      mdr_data_out(32), A2=>mdr_data_out(33));
   ix3739 : nor04 port map ( Y=>nx3738, A0=>mdr_data_out(35), A1=>
      mdr_data_out(34), A2=>mdr_data_out(32), A3=>mdr_data_out(33));
   ix28379 : xnor2 port map ( Y=>nx28378, A0=>nx3776, A1=>nx13023);
   ix3777 : oai22 port map ( Y=>nx3776, A0=>nx28361, A1=>nx28381, B0=>
      nx28390, B1=>nx35387);
   ix28384 : aoi32 port map ( Y=>nx28383, A0=>nx3758, A1=>nx34649, A2=>
      nx28388, B0=>mdr_data_out(36), B1=>nx34643);
   ix3759 : nand02 port map ( Y=>nx3758, A0=>nx28386, A1=>mdr_data_out(36));
   booth_booth_integrtaion_1_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_20, QB=>nx28390, D=>nx16153, 
      CLK=>clk, R=>rst);
   ix16144 : oai21 port map ( Y=>nx16143, A0=>nx28395, A1=>nx35373, B0=>
      nx28397);
   booth_booth_integrtaion_1_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_21, QB=>nx28395, D=>nx16143, 
      CLK=>clk, R=>rst);
   ix28398 : nand03 port map ( Y=>nx28397, A0=>nx35381, A1=>nx4136, A2=>
      nx36077);
   ix4137 : xnor2 port map ( Y=>nx4136, A0=>nx28400, A1=>nx13025);
   ix28401 : aoi22 port map ( Y=>nx28400, A0=>
      booth_booth_integrtaion_1_booth_output_21, A1=>nx3796, B0=>nx3776, B1
      =>nx13023);
   ix28404 : nor02ii port map ( Y=>nx28403, A0=>nx3762, A1=>mdr_data_out(37)
   );
   ix3763 : nor02ii port map ( Y=>nx3762, A0=>mdr_data_out(36), A1=>nx3738);
   ix3787 : nor02ii port map ( Y=>nx3786, A0=>mdr_data_out(37), A1=>nx3762);
   ix28414 : xnor2 port map ( Y=>nx28413, A0=>nx3824, A1=>nx13026);
   ix3825 : oai22 port map ( Y=>nx3824, A0=>nx28400, A1=>nx28416, B0=>
      nx28425, B1=>nx35389);
   ix28419 : aoi32 port map ( Y=>nx28418, A0=>nx3806, A1=>nx34649, A2=>
      nx28423, B0=>mdr_data_out(38), B1=>nx34643);
   ix3807 : nand02 port map ( Y=>nx3806, A0=>nx28421, A1=>mdr_data_out(38));
   booth_booth_integrtaion_1_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_22, QB=>nx28425, D=>nx16133, 
      CLK=>clk, R=>rst);
   ix16124 : oai21 port map ( Y=>nx16123, A0=>nx28430, A1=>nx35373, B0=>
      nx28432);
   booth_booth_integrtaion_1_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_23, QB=>nx28430, D=>nx16123, 
      CLK=>clk, R=>rst);
   ix28433 : nand03 port map ( Y=>nx28432, A0=>nx35381, A1=>nx4112, A2=>
      nx35375);
   ix4113 : xnor2 port map ( Y=>nx4112, A0=>nx28435, A1=>nx13027);
   ix28436 : aoi22 port map ( Y=>nx28435, A0=>
      booth_booth_integrtaion_1_booth_output_23, A1=>nx3844, B0=>nx3824, B1
      =>nx13026);
   ix28439 : nor02ii port map ( Y=>nx28438, A0=>nx3810, A1=>mdr_data_out(39)
   );
   ix3811 : nor02ii port map ( Y=>nx3810, A0=>mdr_data_out(38), A1=>nx3786);
   ix3835 : nor02ii port map ( Y=>nx3834, A0=>mdr_data_out(39), A1=>nx3810);
   ix28449 : xnor2 port map ( Y=>nx28448, A0=>nx3872, A1=>nx13029);
   ix3873 : oai22 port map ( Y=>nx3872, A0=>nx28435, A1=>nx28451, B0=>
      nx28460, B1=>nx35391);
   ix28454 : aoi32 port map ( Y=>nx28453, A0=>nx3854, A1=>nx34649, A2=>
      nx28458, B0=>mdr_data_out(40), B1=>nx34643);
   ix3855 : nand02 port map ( Y=>nx3854, A0=>nx28456, A1=>mdr_data_out(40));
   booth_booth_integrtaion_1_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_24, QB=>nx28460, D=>nx16113, 
      CLK=>clk, R=>rst);
   ix16104 : oai21 port map ( Y=>nx16103, A0=>nx28465, A1=>nx35375, B0=>
      nx28467);
   booth_booth_integrtaion_1_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_25, QB=>nx28465, D=>nx16103, 
      CLK=>clk, R=>rst);
   ix28468 : nand03 port map ( Y=>nx28467, A0=>nx35381, A1=>nx4088, A2=>
      nx35375);
   ix4089 : xnor2 port map ( Y=>nx4088, A0=>nx28470, A1=>nx13031);
   ix28471 : aoi22 port map ( Y=>nx28470, A0=>
      booth_booth_integrtaion_1_booth_output_25, A1=>nx3892, B0=>nx3872, B1
      =>nx13029);
   ix28474 : nor02ii port map ( Y=>nx28473, A0=>nx3858, A1=>mdr_data_out(41)
   );
   ix3859 : nor02ii port map ( Y=>nx3858, A0=>mdr_data_out(40), A1=>nx3834);
   ix3883 : nor02ii port map ( Y=>nx3882, A0=>mdr_data_out(41), A1=>nx3858);
   ix28484 : xnor2 port map ( Y=>nx28483, A0=>nx3920, A1=>nx13033);
   ix3921 : oai22 port map ( Y=>nx3920, A0=>nx28470, A1=>nx28486, B0=>
      nx28495, B1=>nx35393);
   ix28489 : aoi32 port map ( Y=>nx28488, A0=>nx3902, A1=>nx34649, A2=>
      nx28493, B0=>mdr_data_out(42), B1=>nx34643);
   ix3903 : nand02 port map ( Y=>nx3902, A0=>nx28491, A1=>mdr_data_out(42));
   booth_booth_integrtaion_1_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_26, QB=>nx28495, D=>nx16093, 
      CLK=>clk, R=>rst);
   ix16084 : oai21 port map ( Y=>nx16083, A0=>nx28500, A1=>nx35375, B0=>
      nx28502);
   booth_booth_integrtaion_1_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_27, QB=>nx28500, D=>nx16083, 
      CLK=>clk, R=>rst);
   ix28503 : nand03 port map ( Y=>nx28502, A0=>nx35381, A1=>nx4064, A2=>
      nx35375);
   ix4065 : xnor2 port map ( Y=>nx4064, A0=>nx28505, A1=>nx13035);
   ix28506 : aoi22 port map ( Y=>nx28505, A0=>
      booth_booth_integrtaion_1_booth_output_27, A1=>nx3940, B0=>nx3920, B1
      =>nx13033);
   ix28509 : nor02ii port map ( Y=>nx28508, A0=>nx3906, A1=>mdr_data_out(43)
   );
   ix3907 : nor02ii port map ( Y=>nx3906, A0=>mdr_data_out(42), A1=>nx3882);
   ix3931 : nor02ii port map ( Y=>nx3930, A0=>mdr_data_out(43), A1=>nx3906);
   ix28519 : xnor2 port map ( Y=>nx28518, A0=>nx3968, A1=>nx13037);
   ix3969 : oai22 port map ( Y=>nx3968, A0=>nx28505, A1=>nx28521, B0=>
      nx28530, B1=>nx35395);
   ix28524 : aoi32 port map ( Y=>nx28523, A0=>nx3950, A1=>nx34649, A2=>
      nx28528, B0=>mdr_data_out(44), B1=>nx34643);
   ix3951 : nand02 port map ( Y=>nx3950, A0=>nx28526, A1=>mdr_data_out(44));
   booth_booth_integrtaion_1_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_28, QB=>nx28530, D=>nx16073, 
      CLK=>clk, R=>rst);
   ix16064 : oai21 port map ( Y=>nx16063, A0=>nx28535, A1=>nx35375, B0=>
      nx28537);
   booth_booth_integrtaion_1_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_29, QB=>nx28535, D=>nx16063, 
      CLK=>clk, R=>rst);
   ix28538 : nand03 port map ( Y=>nx28537, A0=>nx36085, A1=>nx4040, A2=>
      nx35375);
   ix4041 : xnor2 port map ( Y=>nx4040, A0=>nx28540, A1=>nx13039);
   ix28541 : aoi22 port map ( Y=>nx28540, A0=>
      booth_booth_integrtaion_1_booth_output_29, A1=>nx3988, B0=>nx3968, B1
      =>nx13037);
   ix28544 : nor02ii port map ( Y=>nx28543, A0=>nx3954, A1=>mdr_data_out(45)
   );
   ix3955 : nor02ii port map ( Y=>nx3954, A0=>mdr_data_out(44), A1=>nx3930);
   ix3979 : nor02ii port map ( Y=>nx3978, A0=>mdr_data_out(45), A1=>nx3954);
   ix28554 : xnor2 port map ( Y=>nx28553, A0=>nx4016, A1=>nx4026);
   ix4017 : oai22 port map ( Y=>nx4016, A0=>nx28540, A1=>nx28556, B0=>
      nx28565, B1=>nx35397);
   ix28559 : aoi32 port map ( Y=>nx28558, A0=>nx3998, A1=>nx34651, A2=>
      nx28563, B0=>mdr_data_out(46), B1=>nx34645);
   ix3999 : nand02 port map ( Y=>nx3998, A0=>nx28561, A1=>mdr_data_out(46));
   booth_booth_integrtaion_1_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_31, QB=>nx28565, D=>nx16053, 
      CLK=>clk, R=>rst);
   ix28569 : aoi22 port map ( Y=>nx28568, A0=>mdr_data_out(47), A1=>nx34645, 
      B0=>nx34651, B1=>nx4018);
   ix4019 : xnor2 port map ( Y=>nx4018, A0=>mdr_data_out(47), A1=>nx4002);
   ix4003 : nor02ii port map ( Y=>nx4002, A0=>mdr_data_out(46), A1=>nx3978);
   ix28573 : aoi32 port map ( Y=>nx28572, A0=>nx3974, A1=>nx34651, A2=>
      nx28561, B0=>mdr_data_out(45), B1=>nx34645);
   ix28576 : aoi32 port map ( Y=>nx28575, A0=>nx3926, A1=>nx34651, A2=>
      nx28526, B0=>mdr_data_out(43), B1=>nx34645);
   ix28579 : aoi32 port map ( Y=>nx28578, A0=>nx3878, A1=>nx34651, A2=>
      nx28491, B0=>mdr_data_out(41), B1=>nx34645);
   ix28582 : aoi32 port map ( Y=>nx28581, A0=>nx3830, A1=>nx34651, A2=>
      nx28456, B0=>mdr_data_out(39), B1=>nx34645);
   ix28585 : aoi32 port map ( Y=>nx28584, A0=>nx3782, A1=>nx34651, A2=>
      nx28421, B0=>mdr_data_out(37), B1=>nx34645);
   ix28588 : aoi32 port map ( Y=>nx28587, A0=>nx3734, A1=>nx3670, A2=>
      nx28386, B0=>mdr_data_out(35), B1=>nx34647);
   ix28591 : aoi32 port map ( Y=>nx28590, A0=>nx3684, A1=>nx3670, A2=>
      nx28335, B0=>mdr_data_out(33), B1=>nx34647);
   booth_booth_integrtaion_1_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_1_booth_output_16, QB=>nx28316, D=>nx16193, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_1_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_1_15, QB=>nx28594, D=>nx16203, CLK=>clk, 
      R=>rst);
   ix4409 : aoi21 port map ( Y=>nx4408, A0=>label_2_output(0), A1=>nx35727, 
      B0=>nx36387);
   max_calc_reg_ans2_0 : dff port map ( Q=>max_calc_ans2_0, QB=>OPEN, D=>
      nx25443, CLK=>clk);
   ix24274 : oai21 port map ( Y=>nx24273, A0=>nx28617, A1=>nx34765, B0=>
      nx28619);
   max_calc_reg_comparator_second_inp1_0 : dff port map ( Q=>
      max_calc_comparator_second_inp1_0, QB=>nx28617, D=>nx24273, CLK=>clk);
   ix28620 : nand03 port map ( Y=>nx28619, A0=>nx36389, A1=>nx16932, A2=>
      nx34783);
   labelsregfile_label3_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_3_output(0), QB=>OPEN, D=>nx15523, CLK=>clk, R=>rst);
   lat_label_3_input_0 : latch port map ( Q=>label_3_input_0, D=>nx3082, CLK
      =>nx34519);
   ix3083 : oai21 port map ( Y=>nx3082, A0=>nx28626, A1=>nx34419, B0=>
      nx28630);
   reg_label_3_input_state_machine_0 : dffr port map ( Q=>
      label_3_input_state_machine_0, QB=>nx28626, D=>nx15513, CLK=>clk, R=>
      rst);
   ix28631 : oai21 port map ( Y=>nx28630, A0=>nx35723, A1=>label_3_output(0), 
      B0=>nx3070);
   booth_booth_integrtaion_2_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_1, QB=>OPEN, D=>nx15493, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_2, QB=>nx29051, D=>nx15483, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_3, QB=>OPEN, D=>nx15473, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_4, QB=>nx29049, D=>nx15463, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_5, QB=>OPEN, D=>nx15453, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_6, QB=>nx29047, D=>nx15443, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_7, QB=>OPEN, D=>nx15433, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_8, QB=>nx29045, D=>nx15423, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_9, QB=>OPEN, D=>nx15413, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_10, QB=>nx29043, D=>nx15403, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_11, QB=>OPEN, D=>nx15393, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_12, QB=>nx29041, D=>nx15383, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_13, QB=>OPEN, D=>nx15373, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_14, QB=>nx29039, D=>nx15363, CLK=>clk, 
      R=>rst);
   ix28680 : aoi22 port map ( Y=>nx28679, A0=>mdr_data_out(15), A1=>nx34603, 
      B0=>nx2868, B1=>nx2874);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_reg_output_0, QB=>OPEN, 
      D=>nx15003, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_0, QB=>OPEN, D=>nx14989, CLK
      =>clk, S=>nx34477);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_reg_output_9, QB=>OPEN, 
      D=>nx15183, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_9, QB=>OPEN, D=>nx15173, CLK
      =>clk, R=>nx34477);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_8, QB=>OPEN, 
      D=>nx15163, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_8, QB=>OPEN, D=>nx15153, CLK
      =>clk, R=>nx34477);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_7, QB=>OPEN, 
      D=>nx15143, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_7, QB=>OPEN, D=>nx15133, CLK
      =>clk, R=>nx34477);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_6, QB=>OPEN, 
      D=>nx15123, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_6, QB=>OPEN, D=>nx15113, CLK
      =>clk, R=>nx34477);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_5, QB=>OPEN, 
      D=>nx15103, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_5, QB=>OPEN, D=>nx15093, CLK
      =>clk, R=>nx34475);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_4, QB=>OPEN, 
      D=>nx15083, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_4, QB=>OPEN, D=>nx15073, CLK
      =>clk, R=>nx34475);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_3, QB=>OPEN, 
      D=>nx15063, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_3, QB=>OPEN, D=>nx15053, CLK
      =>clk, R=>nx34475);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_2, QB=>OPEN, 
      D=>nx15043, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_2, QB=>OPEN, D=>nx15033, CLK
      =>clk, R=>nx34475);
   booth_booth_integrtaion_2_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_2_shift_Reg_output_1, QB=>OPEN, 
      D=>nx15023, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_2_shift_Reg_count_1, QB=>OPEN, D=>nx15013, CLK
      =>clk, R=>nx34475);
   ix14984 : nand02 port map ( Y=>nx14983, A0=>nx35819, A1=>nx34589);
   booth_booth_integrtaion_2_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx28726, D=>nx14983, CLK=>clk, S=>nx34475);
   ix2869 : nand02 port map ( Y=>nx2868, A0=>nx28747, A1=>nx28759);
   ix28748 : oai21 port map ( Y=>nx28747, A0=>nx34617, A1=>nx34611, B0=>
      mdr_data_out(48));
   ix15194 : oai21 port map ( Y=>nx15193, A0=>nx28752, A1=>nx35399, B0=>
      nx28754);
   booth_booth_integrtaion_2_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx28752, D=>nx15193, CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx28756, D=>nx15503, CLK=>clk, R=>rst);
   ix28764 : xnor2 port map ( Y=>nx28763, A0=>nx2338, A1=>nx12965);
   ix15334 : oai21 port map ( Y=>nx15333, A0=>nx28769, A1=>nx35399, B0=>
      nx28771);
   booth_booth_integrtaion_2_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_17, QB=>nx28769, D=>nx15333, 
      CLK=>clk, R=>rst);
   ix28772 : nand03 port map ( Y=>nx28771, A0=>nx35407, A1=>nx2846, A2=>
      nx36093);
   ix2847 : xnor2 port map ( Y=>nx2846, A0=>nx28774, A1=>nx12967);
   ix28775 : aoi22 port map ( Y=>nx28774, A0=>
      booth_booth_integrtaion_2_booth_output_17, A1=>nx2362, B0=>nx2338, B1
      =>nx12965);
   ix2347 : nand02 port map ( Y=>nx2346, A0=>mdr_data_out(49), A1=>
      mdr_data_out(48));
   ix28779 : or02 port map ( Y=>nx28778, A0=>mdr_data_out(48), A1=>
      mdr_data_out(49));
   ix28785 : xnor2 port map ( Y=>nx28784, A0=>nx2390, A1=>nx12969);
   ix2391 : oai22 port map ( Y=>nx2390, A0=>nx28774, A1=>nx28787, B0=>
      nx28794, B1=>nx35411);
   ix28790 : aoi32 port map ( Y=>nx28789, A0=>nx2372, A1=>nx34617, A2=>
      nx28792, B0=>mdr_data_out(50), B1=>nx34611);
   ix2373 : oai21 port map ( Y=>nx2372, A0=>mdr_data_out(48), A1=>
      mdr_data_out(49), B0=>mdr_data_out(50));
   booth_booth_integrtaion_2_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_18, QB=>nx28794, D=>nx15323, 
      CLK=>clk, R=>rst);
   ix15314 : oai21 port map ( Y=>nx15313, A0=>nx28799, A1=>nx35399, B0=>
      nx28801);
   booth_booth_integrtaion_2_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_19, QB=>nx28799, D=>nx15313, 
      CLK=>clk, R=>rst);
   ix28802 : nand03 port map ( Y=>nx28801, A0=>nx35407, A1=>nx2822, A2=>
      nx36093);
   ix2823 : xnor2 port map ( Y=>nx2822, A0=>nx28804, A1=>nx12970);
   ix28805 : aoi22 port map ( Y=>nx28804, A0=>
      booth_booth_integrtaion_2_booth_output_19, A1=>nx2410, B0=>nx2390, B1
      =>nx12969);
   ix28808 : nor02ii port map ( Y=>nx28807, A0=>nx2376, A1=>mdr_data_out(51)
   );
   ix2377 : nor03_2x port map ( Y=>nx2376, A0=>mdr_data_out(50), A1=>
      mdr_data_out(48), A2=>mdr_data_out(49));
   ix2401 : nor04 port map ( Y=>nx2400, A0=>mdr_data_out(51), A1=>
      mdr_data_out(50), A2=>mdr_data_out(48), A3=>mdr_data_out(49));
   ix28822 : xnor2 port map ( Y=>nx28821, A0=>nx2438, A1=>nx12971);
   ix2439 : oai22 port map ( Y=>nx2438, A0=>nx28804, A1=>nx28824, B0=>
      nx28833, B1=>nx35413);
   ix28827 : aoi32 port map ( Y=>nx28826, A0=>nx2420, A1=>nx34617, A2=>
      nx28831, B0=>mdr_data_out(52), B1=>nx34611);
   ix2421 : nand02 port map ( Y=>nx2420, A0=>nx28829, A1=>mdr_data_out(52));
   booth_booth_integrtaion_2_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_20, QB=>nx28833, D=>nx15303, 
      CLK=>clk, R=>rst);
   ix15294 : oai21 port map ( Y=>nx15293, A0=>nx28838, A1=>nx35399, B0=>
      nx28840);
   booth_booth_integrtaion_2_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_21, QB=>nx28838, D=>nx15293, 
      CLK=>clk, R=>rst);
   ix28841 : nand03 port map ( Y=>nx28840, A0=>nx35407, A1=>nx2798, A2=>
      nx36093);
   ix2799 : xnor2 port map ( Y=>nx2798, A0=>nx28843, A1=>nx12973);
   ix28844 : aoi22 port map ( Y=>nx28843, A0=>
      booth_booth_integrtaion_2_booth_output_21, A1=>nx2458, B0=>nx2438, B1
      =>nx12971);
   ix28847 : nor02ii port map ( Y=>nx28846, A0=>nx2424, A1=>mdr_data_out(53)
   );
   ix2425 : nor02ii port map ( Y=>nx2424, A0=>mdr_data_out(52), A1=>nx2400);
   ix2449 : nor02ii port map ( Y=>nx2448, A0=>mdr_data_out(53), A1=>nx2424);
   ix28857 : xnor2 port map ( Y=>nx28856, A0=>nx2486, A1=>nx12975);
   ix2487 : oai22 port map ( Y=>nx2486, A0=>nx28843, A1=>nx28859, B0=>
      nx28868, B1=>nx35415);
   ix28862 : aoi32 port map ( Y=>nx28861, A0=>nx2468, A1=>nx34617, A2=>
      nx28866, B0=>mdr_data_out(54), B1=>nx34611);
   ix2469 : nand02 port map ( Y=>nx2468, A0=>nx28864, A1=>mdr_data_out(54));
   booth_booth_integrtaion_2_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_22, QB=>nx28868, D=>nx15283, 
      CLK=>clk, R=>rst);
   ix15274 : oai21 port map ( Y=>nx15273, A0=>nx28873, A1=>nx35399, B0=>
      nx28875);
   booth_booth_integrtaion_2_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_23, QB=>nx28873, D=>nx15273, 
      CLK=>clk, R=>rst);
   ix28876 : nand03 port map ( Y=>nx28875, A0=>nx35407, A1=>nx2774, A2=>
      nx35401);
   ix2775 : xnor2 port map ( Y=>nx2774, A0=>nx28878, A1=>nx12977);
   ix28879 : aoi22 port map ( Y=>nx28878, A0=>
      booth_booth_integrtaion_2_booth_output_23, A1=>nx2506, B0=>nx2486, B1
      =>nx12975);
   ix28882 : nor02ii port map ( Y=>nx28881, A0=>nx2472, A1=>mdr_data_out(55)
   );
   ix2473 : nor02ii port map ( Y=>nx2472, A0=>mdr_data_out(54), A1=>nx2448);
   ix2497 : nor02ii port map ( Y=>nx2496, A0=>mdr_data_out(55), A1=>nx2472);
   ix28892 : xnor2 port map ( Y=>nx28891, A0=>nx2534, A1=>nx12978);
   ix2535 : oai22 port map ( Y=>nx2534, A0=>nx28878, A1=>nx28894, B0=>
      nx28903, B1=>nx35417);
   ix28897 : aoi32 port map ( Y=>nx28896, A0=>nx2516, A1=>nx34617, A2=>
      nx28901, B0=>mdr_data_out(56), B1=>nx34611);
   ix2517 : nand02 port map ( Y=>nx2516, A0=>nx28899, A1=>mdr_data_out(56));
   booth_booth_integrtaion_2_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_24, QB=>nx28903, D=>nx15263, 
      CLK=>clk, R=>rst);
   ix15254 : oai21 port map ( Y=>nx15253, A0=>nx28908, A1=>nx35401, B0=>
      nx28910);
   booth_booth_integrtaion_2_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_25, QB=>nx28908, D=>nx15253, 
      CLK=>clk, R=>rst);
   ix28911 : nand03 port map ( Y=>nx28910, A0=>nx35407, A1=>nx2750, A2=>
      nx35401);
   ix2751 : xnor2 port map ( Y=>nx2750, A0=>nx28913, A1=>nx12979);
   ix28914 : aoi22 port map ( Y=>nx28913, A0=>
      booth_booth_integrtaion_2_booth_output_25, A1=>nx2554, B0=>nx2534, B1
      =>nx12978);
   ix28917 : nor02ii port map ( Y=>nx28916, A0=>nx2520, A1=>mdr_data_out(57)
   );
   ix2521 : nor02ii port map ( Y=>nx2520, A0=>mdr_data_out(56), A1=>nx2496);
   ix2545 : nor02ii port map ( Y=>nx2544, A0=>mdr_data_out(57), A1=>nx2520);
   ix28927 : xnor2 port map ( Y=>nx28926, A0=>nx2582, A1=>nx12981);
   ix2583 : oai22 port map ( Y=>nx2582, A0=>nx28913, A1=>nx28929, B0=>
      nx28938, B1=>nx35419);
   ix28932 : aoi32 port map ( Y=>nx28931, A0=>nx2564, A1=>nx34617, A2=>
      nx28936, B0=>mdr_data_out(58), B1=>nx34611);
   ix2565 : nand02 port map ( Y=>nx2564, A0=>nx28934, A1=>mdr_data_out(58));
   booth_booth_integrtaion_2_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_26, QB=>nx28938, D=>nx15243, 
      CLK=>clk, R=>rst);
   ix15234 : oai21 port map ( Y=>nx15233, A0=>nx28943, A1=>nx35401, B0=>
      nx28945);
   booth_booth_integrtaion_2_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_27, QB=>nx28943, D=>nx15233, 
      CLK=>clk, R=>rst);
   ix28946 : nand03 port map ( Y=>nx28945, A0=>nx35407, A1=>nx2726, A2=>
      nx35401);
   ix2727 : xnor2 port map ( Y=>nx2726, A0=>nx28948, A1=>nx12983);
   ix28949 : aoi22 port map ( Y=>nx28948, A0=>
      booth_booth_integrtaion_2_booth_output_27, A1=>nx2602, B0=>nx2582, B1
      =>nx12981);
   ix28952 : nor02ii port map ( Y=>nx28951, A0=>nx2568, A1=>mdr_data_out(59)
   );
   ix2569 : nor02ii port map ( Y=>nx2568, A0=>mdr_data_out(58), A1=>nx2544);
   ix2593 : nor02ii port map ( Y=>nx2592, A0=>mdr_data_out(59), A1=>nx2568);
   ix28962 : xnor2 port map ( Y=>nx28961, A0=>nx2630, A1=>nx12985);
   ix2631 : oai22 port map ( Y=>nx2630, A0=>nx28948, A1=>nx28964, B0=>
      nx28973, B1=>nx35421);
   ix28967 : aoi32 port map ( Y=>nx28966, A0=>nx2612, A1=>nx34617, A2=>
      nx28971, B0=>mdr_data_out(60), B1=>nx34611);
   ix2613 : nand02 port map ( Y=>nx2612, A0=>nx28969, A1=>mdr_data_out(60));
   booth_booth_integrtaion_2_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_28, QB=>nx28973, D=>nx15223, 
      CLK=>clk, R=>rst);
   ix15214 : oai21 port map ( Y=>nx15213, A0=>nx28978, A1=>nx35401, B0=>
      nx28980);
   booth_booth_integrtaion_2_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_29, QB=>nx28978, D=>nx15213, 
      CLK=>clk, R=>rst);
   ix28981 : nand03 port map ( Y=>nx28980, A0=>nx36101, A1=>nx2702, A2=>
      nx35401);
   ix2703 : xnor2 port map ( Y=>nx2702, A0=>nx28983, A1=>nx12987);
   ix28984 : aoi22 port map ( Y=>nx28983, A0=>
      booth_booth_integrtaion_2_booth_output_29, A1=>nx2650, B0=>nx2630, B1
      =>nx12985);
   ix28987 : nor02ii port map ( Y=>nx28986, A0=>nx2616, A1=>mdr_data_out(61)
   );
   ix2617 : nor02ii port map ( Y=>nx2616, A0=>mdr_data_out(60), A1=>nx2592);
   ix2641 : nor02ii port map ( Y=>nx2640, A0=>mdr_data_out(61), A1=>nx2616);
   ix28997 : xnor2 port map ( Y=>nx28996, A0=>nx2678, A1=>nx2688);
   ix2679 : oai22 port map ( Y=>nx2678, A0=>nx28983, A1=>nx28999, B0=>
      nx29008, B1=>nx35423);
   ix29002 : aoi32 port map ( Y=>nx29001, A0=>nx2660, A1=>nx34619, A2=>
      nx29006, B0=>mdr_data_out(62), B1=>nx34613);
   ix2661 : nand02 port map ( Y=>nx2660, A0=>nx29004, A1=>mdr_data_out(62));
   booth_booth_integrtaion_2_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_31, QB=>nx29008, D=>nx15203, 
      CLK=>clk, R=>rst);
   ix29012 : aoi22 port map ( Y=>nx29011, A0=>mdr_data_out(63), A1=>nx34613, 
      B0=>nx34619, B1=>nx2680);
   ix2681 : xnor2 port map ( Y=>nx2680, A0=>mdr_data_out(63), A1=>nx2664);
   ix2665 : nor02ii port map ( Y=>nx2664, A0=>mdr_data_out(62), A1=>nx2640);
   ix29016 : aoi32 port map ( Y=>nx29015, A0=>nx2636, A1=>nx34619, A2=>
      nx29004, B0=>mdr_data_out(61), B1=>nx34613);
   ix29019 : aoi32 port map ( Y=>nx29018, A0=>nx2588, A1=>nx34619, A2=>
      nx28969, B0=>mdr_data_out(59), B1=>nx34613);
   ix29022 : aoi32 port map ( Y=>nx29021, A0=>nx2540, A1=>nx34619, A2=>
      nx28934, B0=>mdr_data_out(57), B1=>nx34613);
   ix29025 : aoi32 port map ( Y=>nx29024, A0=>nx2492, A1=>nx34619, A2=>
      nx28899, B0=>mdr_data_out(55), B1=>nx34613);
   ix29028 : aoi32 port map ( Y=>nx29027, A0=>nx2444, A1=>nx34619, A2=>
      nx28864, B0=>mdr_data_out(53), B1=>nx34613);
   ix29031 : aoi32 port map ( Y=>nx29030, A0=>nx2396, A1=>nx2332, A2=>
      nx28829, B0=>mdr_data_out(51), B1=>nx34615);
   ix29034 : aoi32 port map ( Y=>nx29033, A0=>nx2346, A1=>nx2332, A2=>
      nx28778, B0=>mdr_data_out(49), B1=>nx34615);
   booth_booth_integrtaion_2_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_2_booth_output_16, QB=>nx28759, D=>nx15343, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_2_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_2_15, QB=>nx29037, D=>nx15353, CLK=>clk, 
      R=>rst);
   ix3071 : aoi21 port map ( Y=>nx3070, A0=>label_3_output(0), A1=>nx35723, 
      B0=>nx36387);
   ix21594 : oai21 port map ( Y=>nx21593, A0=>nx29061, A1=>nx34765, B0=>
      nx29063);
   max_calc_reg_comparator_third_inp1_0 : dff port map ( Q=>
      max_calc_comparator_third_inp1_0, QB=>nx29061, D=>nx21593, CLK=>clk);
   ix29064 : nand03 port map ( Y=>nx29063, A0=>label_5_output(0), A1=>
      nx35453, A2=>nx34765);
   labelsregfile_label5_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_5_output(0), QB=>OPEN, D=>nx20193, CLK=>clk, R=>rst);
   lat_label_5_input_0 : latch port map ( Q=>label_5_input_0, D=>nx10396, 
      CLK=>nx34521);
   ix10397 : oai21 port map ( Y=>nx10396, A0=>nx29069, A1=>nx34419, B0=>
      nx29073);
   reg_label_5_input_state_machine_0 : dffr port map ( Q=>
      label_5_input_state_machine_0, QB=>nx29069, D=>nx20183, CLK=>clk, R=>
      rst);
   ix29074 : oai21 port map ( Y=>nx29073, A0=>nx35763, A1=>label_5_output(0), 
      B0=>nx10384);
   booth_booth_integrtaion_4_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_1, QB=>OPEN, D=>nx20163, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_2, QB=>nx29494, D=>nx20153, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_3, QB=>OPEN, D=>nx20143, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_4, QB=>nx29492, D=>nx20133, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_5, QB=>OPEN, D=>nx20123, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_6, QB=>nx29490, D=>nx20113, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_7, QB=>OPEN, D=>nx20103, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_8, QB=>nx29488, D=>nx20093, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_9, QB=>OPEN, D=>nx20083, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_10, QB=>nx29486, D=>nx20073, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_11, QB=>OPEN, D=>nx20063, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_12, QB=>nx29484, D=>nx20053, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_13, QB=>OPEN, D=>nx20043, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_14, QB=>nx29482, D=>nx20033, CLK=>clk, 
      R=>rst);
   ix29123 : aoi22 port map ( Y=>nx29122, A0=>mdr_data_out(15), A1=>nx34939, 
      B0=>nx10182, B1=>nx10188);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_reg_output_0, QB=>OPEN, 
      D=>nx19673, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_0, QB=>OPEN, D=>nx19659, CLK
      =>clk, S=>nx34481);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_reg_output_9, QB=>OPEN, 
      D=>nx19853, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_9, QB=>OPEN, D=>nx19843, CLK
      =>clk, R=>nx34481);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_8, QB=>OPEN, 
      D=>nx19833, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_8, QB=>OPEN, D=>nx19823, CLK
      =>clk, R=>nx34479);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_7, QB=>OPEN, 
      D=>nx19813, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_7, QB=>OPEN, D=>nx19803, CLK
      =>clk, R=>nx34479);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_6, QB=>OPEN, 
      D=>nx19793, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_6, QB=>OPEN, D=>nx19783, CLK
      =>clk, R=>nx34479);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_5, QB=>OPEN, 
      D=>nx19773, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_5, QB=>OPEN, D=>nx19763, CLK
      =>clk, R=>nx34479);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_4, QB=>OPEN, 
      D=>nx19753, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_4, QB=>OPEN, D=>nx19743, CLK
      =>clk, R=>nx34479);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_3, QB=>OPEN, 
      D=>nx19733, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_3, QB=>OPEN, D=>nx19723, CLK
      =>clk, R=>nx34479);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_2, QB=>OPEN, 
      D=>nx19713, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_2, QB=>OPEN, D=>nx19703, CLK
      =>clk, R=>nx34479);
   booth_booth_integrtaion_4_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_4_shift_Reg_output_1, QB=>OPEN, 
      D=>nx19693, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_4_shift_Reg_count_1, QB=>OPEN, D=>nx19683, CLK
      =>clk, R=>nx34477);
   ix19654 : nand02 port map ( Y=>nx19653, A0=>nx35823, A1=>nx34925);
   booth_booth_integrtaion_4_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx29169, D=>nx19653, CLK=>clk, S=>nx34477);
   ix10183 : nand02 port map ( Y=>nx10182, A0=>nx29190, A1=>nx29202);
   ix29191 : oai21 port map ( Y=>nx29190, A0=>nx34953, A1=>nx34947, B0=>
      mdr_data_out(80));
   ix19864 : oai21 port map ( Y=>nx19863, A0=>nx29195, A1=>nx35425, B0=>
      nx29197);
   booth_booth_integrtaion_4_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx29195, D=>nx19863, CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx29199, D=>nx20173, CLK=>clk, R=>rst);
   ix29207 : xnor2 port map ( Y=>nx29206, A0=>nx9652, A1=>nx13217);
   ix20004 : oai21 port map ( Y=>nx20003, A0=>nx29212, A1=>nx35425, B0=>
      nx29214);
   booth_booth_integrtaion_4_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_17, QB=>nx29212, D=>nx20003, 
      CLK=>clk, R=>rst);
   ix29215 : nand03 port map ( Y=>nx29214, A0=>nx35433, A1=>nx10160, A2=>
      nx36109);
   ix10161 : xnor2 port map ( Y=>nx10160, A0=>nx29217, A1=>nx13219);
   ix29218 : aoi22 port map ( Y=>nx29217, A0=>
      booth_booth_integrtaion_4_booth_output_17, A1=>nx9676, B0=>nx9652, B1
      =>nx13217);
   ix9661 : nand02 port map ( Y=>nx9660, A0=>mdr_data_out(81), A1=>
      mdr_data_out(80));
   ix29222 : or02 port map ( Y=>nx29221, A0=>mdr_data_out(80), A1=>
      mdr_data_out(81));
   ix29228 : xnor2 port map ( Y=>nx29227, A0=>nx9704, A1=>nx13221);
   ix9705 : oai22 port map ( Y=>nx9704, A0=>nx29217, A1=>nx29230, B0=>
      nx29237, B1=>nx35437);
   ix29233 : aoi32 port map ( Y=>nx29232, A0=>nx9686, A1=>nx34953, A2=>
      nx29235, B0=>mdr_data_out(82), B1=>nx34947);
   ix9687 : oai21 port map ( Y=>nx9686, A0=>mdr_data_out(80), A1=>
      mdr_data_out(81), B0=>mdr_data_out(82));
   booth_booth_integrtaion_4_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_18, QB=>nx29237, D=>nx19993, 
      CLK=>clk, R=>rst);
   ix19984 : oai21 port map ( Y=>nx19983, A0=>nx29242, A1=>nx35425, B0=>
      nx29244);
   booth_booth_integrtaion_4_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_19, QB=>nx29242, D=>nx19983, 
      CLK=>clk, R=>rst);
   ix29245 : nand03 port map ( Y=>nx29244, A0=>nx35433, A1=>nx10136, A2=>
      nx36109);
   ix10137 : xnor2 port map ( Y=>nx10136, A0=>nx29247, A1=>nx13223);
   ix29248 : aoi22 port map ( Y=>nx29247, A0=>
      booth_booth_integrtaion_4_booth_output_19, A1=>nx9724, B0=>nx9704, B1
      =>nx13221);
   ix29251 : nor02ii port map ( Y=>nx29250, A0=>nx9690, A1=>mdr_data_out(83)
   );
   ix9691 : nor03_2x port map ( Y=>nx9690, A0=>mdr_data_out(82), A1=>
      mdr_data_out(80), A2=>mdr_data_out(81));
   ix9715 : nor04 port map ( Y=>nx9714, A0=>mdr_data_out(83), A1=>
      mdr_data_out(82), A2=>mdr_data_out(80), A3=>mdr_data_out(81));
   ix29265 : xnor2 port map ( Y=>nx29264, A0=>nx9752, A1=>nx13224);
   ix9753 : oai22 port map ( Y=>nx9752, A0=>nx29247, A1=>nx29267, B0=>
      nx29276, B1=>nx35439);
   ix29270 : aoi32 port map ( Y=>nx29269, A0=>nx9734, A1=>nx34953, A2=>
      nx29274, B0=>mdr_data_out(84), B1=>nx34947);
   ix9735 : nand02 port map ( Y=>nx9734, A0=>nx29272, A1=>mdr_data_out(84));
   booth_booth_integrtaion_4_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_20, QB=>nx29276, D=>nx19973, 
      CLK=>clk, R=>rst);
   ix19964 : oai21 port map ( Y=>nx19963, A0=>nx29281, A1=>nx35425, B0=>
      nx29283);
   booth_booth_integrtaion_4_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_21, QB=>nx29281, D=>nx19963, 
      CLK=>clk, R=>rst);
   ix29284 : nand03 port map ( Y=>nx29283, A0=>nx35433, A1=>nx10112, A2=>
      nx36109);
   ix10113 : xnor2 port map ( Y=>nx10112, A0=>nx29286, A1=>nx13225);
   ix29287 : aoi22 port map ( Y=>nx29286, A0=>
      booth_booth_integrtaion_4_booth_output_21, A1=>nx9772, B0=>nx9752, B1
      =>nx13224);
   ix29290 : nor02ii port map ( Y=>nx29289, A0=>nx9738, A1=>mdr_data_out(85)
   );
   ix9739 : nor02ii port map ( Y=>nx9738, A0=>mdr_data_out(84), A1=>nx9714);
   ix9763 : nor02ii port map ( Y=>nx9762, A0=>mdr_data_out(85), A1=>nx9738);
   ix29300 : xnor2 port map ( Y=>nx29299, A0=>nx9800, A1=>nx13226);
   ix9801 : oai22 port map ( Y=>nx9800, A0=>nx29286, A1=>nx29302, B0=>
      nx29311, B1=>nx35441);
   ix29305 : aoi32 port map ( Y=>nx29304, A0=>nx9782, A1=>nx34953, A2=>
      nx29309, B0=>mdr_data_out(86), B1=>nx34947);
   ix9783 : nand02 port map ( Y=>nx9782, A0=>nx29307, A1=>mdr_data_out(86));
   booth_booth_integrtaion_4_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_22, QB=>nx29311, D=>nx19953, 
      CLK=>clk, R=>rst);
   ix19944 : oai21 port map ( Y=>nx19943, A0=>nx29316, A1=>nx35425, B0=>
      nx29318);
   booth_booth_integrtaion_4_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_23, QB=>nx29316, D=>nx19943, 
      CLK=>clk, R=>rst);
   ix29319 : nand03 port map ( Y=>nx29318, A0=>nx35433, A1=>nx10088, A2=>
      nx35427);
   ix10089 : xnor2 port map ( Y=>nx10088, A0=>nx29321, A1=>nx13227);
   ix29322 : aoi22 port map ( Y=>nx29321, A0=>
      booth_booth_integrtaion_4_booth_output_23, A1=>nx9820, B0=>nx9800, B1
      =>nx13226);
   ix29325 : nor02ii port map ( Y=>nx29324, A0=>nx9786, A1=>mdr_data_out(87)
   );
   ix9787 : nor02ii port map ( Y=>nx9786, A0=>mdr_data_out(86), A1=>nx9762);
   ix9811 : nor02ii port map ( Y=>nx9810, A0=>mdr_data_out(87), A1=>nx9786);
   ix29335 : xnor2 port map ( Y=>nx29334, A0=>nx9848, A1=>nx13228);
   ix9849 : oai22 port map ( Y=>nx9848, A0=>nx29321, A1=>nx29337, B0=>
      nx29346, B1=>nx35443);
   ix29340 : aoi32 port map ( Y=>nx29339, A0=>nx9830, A1=>nx34953, A2=>
      nx29344, B0=>mdr_data_out(88), B1=>nx34947);
   ix9831 : nand02 port map ( Y=>nx9830, A0=>nx29342, A1=>mdr_data_out(88));
   booth_booth_integrtaion_4_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_24, QB=>nx29346, D=>nx19933, 
      CLK=>clk, R=>rst);
   ix19924 : oai21 port map ( Y=>nx19923, A0=>nx29351, A1=>nx35427, B0=>
      nx29353);
   booth_booth_integrtaion_4_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_25, QB=>nx29351, D=>nx19923, 
      CLK=>clk, R=>rst);
   ix29354 : nand03 port map ( Y=>nx29353, A0=>nx35433, A1=>nx10064, A2=>
      nx35427);
   ix10065 : xnor2 port map ( Y=>nx10064, A0=>nx29356, A1=>nx13229);
   ix29357 : aoi22 port map ( Y=>nx29356, A0=>
      booth_booth_integrtaion_4_booth_output_25, A1=>nx9868, B0=>nx9848, B1
      =>nx13228);
   ix29360 : nor02ii port map ( Y=>nx29359, A0=>nx9834, A1=>mdr_data_out(89)
   );
   ix9835 : nor02ii port map ( Y=>nx9834, A0=>mdr_data_out(88), A1=>nx9810);
   ix9859 : nor02ii port map ( Y=>nx9858, A0=>mdr_data_out(89), A1=>nx9834);
   ix29370 : xnor2 port map ( Y=>nx29369, A0=>nx9896, A1=>nx13231);
   ix9897 : oai22 port map ( Y=>nx9896, A0=>nx29356, A1=>nx29372, B0=>
      nx29381, B1=>nx35445);
   ix29375 : aoi32 port map ( Y=>nx29374, A0=>nx9878, A1=>nx34953, A2=>
      nx29379, B0=>mdr_data_out(90), B1=>nx34947);
   ix9879 : nand02 port map ( Y=>nx9878, A0=>nx29377, A1=>mdr_data_out(90));
   booth_booth_integrtaion_4_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_26, QB=>nx29381, D=>nx19913, 
      CLK=>clk, R=>rst);
   ix19904 : oai21 port map ( Y=>nx19903, A0=>nx29386, A1=>nx35427, B0=>
      nx29388);
   booth_booth_integrtaion_4_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_27, QB=>nx29386, D=>nx19903, 
      CLK=>clk, R=>rst);
   ix29389 : nand03 port map ( Y=>nx29388, A0=>nx35433, A1=>nx10040, A2=>
      nx35427);
   ix10041 : xnor2 port map ( Y=>nx10040, A0=>nx29391, A1=>nx13233);
   ix29392 : aoi22 port map ( Y=>nx29391, A0=>
      booth_booth_integrtaion_4_booth_output_27, A1=>nx9916, B0=>nx9896, B1
      =>nx13231);
   ix29395 : nor02ii port map ( Y=>nx29394, A0=>nx9882, A1=>mdr_data_out(91)
   );
   ix9883 : nor02ii port map ( Y=>nx9882, A0=>mdr_data_out(90), A1=>nx9858);
   ix9907 : nor02ii port map ( Y=>nx9906, A0=>mdr_data_out(91), A1=>nx9882);
   ix29405 : xnor2 port map ( Y=>nx29404, A0=>nx9944, A1=>nx13235);
   ix9945 : oai22 port map ( Y=>nx9944, A0=>nx29391, A1=>nx29407, B0=>
      nx29416, B1=>nx35447);
   ix29410 : aoi32 port map ( Y=>nx29409, A0=>nx9926, A1=>nx34953, A2=>
      nx29414, B0=>mdr_data_out(92), B1=>nx34947);
   ix9927 : nand02 port map ( Y=>nx9926, A0=>nx29412, A1=>mdr_data_out(92));
   booth_booth_integrtaion_4_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_28, QB=>nx29416, D=>nx19893, 
      CLK=>clk, R=>rst);
   ix19884 : oai21 port map ( Y=>nx19883, A0=>nx29421, A1=>nx35427, B0=>
      nx29423);
   booth_booth_integrtaion_4_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_29, QB=>nx29421, D=>nx19883, 
      CLK=>clk, R=>rst);
   ix29424 : nand03 port map ( Y=>nx29423, A0=>nx36117, A1=>nx10016, A2=>
      nx35427);
   ix10017 : xnor2 port map ( Y=>nx10016, A0=>nx29426, A1=>nx13236);
   ix29427 : aoi22 port map ( Y=>nx29426, A0=>
      booth_booth_integrtaion_4_booth_output_29, A1=>nx9964, B0=>nx9944, B1
      =>nx13235);
   ix29430 : nor02ii port map ( Y=>nx29429, A0=>nx9930, A1=>mdr_data_out(93)
   );
   ix9931 : nor02ii port map ( Y=>nx9930, A0=>mdr_data_out(92), A1=>nx9906);
   ix9955 : nor02ii port map ( Y=>nx9954, A0=>mdr_data_out(93), A1=>nx9930);
   ix29440 : xnor2 port map ( Y=>nx29439, A0=>nx9992, A1=>nx10002);
   ix9993 : oai22 port map ( Y=>nx9992, A0=>nx29426, A1=>nx29442, B0=>
      nx29451, B1=>nx35449);
   ix29445 : aoi32 port map ( Y=>nx29444, A0=>nx9974, A1=>nx34955, A2=>
      nx29449, B0=>mdr_data_out(94), B1=>nx34949);
   ix9975 : nand02 port map ( Y=>nx9974, A0=>nx29447, A1=>mdr_data_out(94));
   booth_booth_integrtaion_4_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_31, QB=>nx29451, D=>nx19873, 
      CLK=>clk, R=>rst);
   ix29455 : aoi22 port map ( Y=>nx29454, A0=>mdr_data_out(95), A1=>nx34949, 
      B0=>nx34955, B1=>nx9994);
   ix9995 : xnor2 port map ( Y=>nx9994, A0=>mdr_data_out(95), A1=>nx9978);
   ix9979 : nor02ii port map ( Y=>nx9978, A0=>mdr_data_out(94), A1=>nx9954);
   ix29459 : aoi32 port map ( Y=>nx29458, A0=>nx9950, A1=>nx34955, A2=>
      nx29447, B0=>mdr_data_out(93), B1=>nx34949);
   ix29462 : aoi32 port map ( Y=>nx29461, A0=>nx9902, A1=>nx34955, A2=>
      nx29412, B0=>mdr_data_out(91), B1=>nx34949);
   ix29465 : aoi32 port map ( Y=>nx29464, A0=>nx9854, A1=>nx34955, A2=>
      nx29377, B0=>mdr_data_out(89), B1=>nx34949);
   ix29468 : aoi32 port map ( Y=>nx29467, A0=>nx9806, A1=>nx34955, A2=>
      nx29342, B0=>mdr_data_out(87), B1=>nx34949);
   ix29471 : aoi32 port map ( Y=>nx29470, A0=>nx9758, A1=>nx34955, A2=>
      nx29307, B0=>mdr_data_out(85), B1=>nx34949);
   ix29474 : aoi32 port map ( Y=>nx29473, A0=>nx9710, A1=>nx9646, A2=>
      nx29272, B0=>mdr_data_out(83), B1=>nx34951);
   ix29477 : aoi32 port map ( Y=>nx29476, A0=>nx9660, A1=>nx9646, A2=>
      nx29221, B0=>mdr_data_out(81), B1=>nx34951);
   booth_booth_integrtaion_4_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_4_booth_output_16, QB=>nx29202, D=>nx20013, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_4_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_4_15, QB=>nx29480, D=>nx20023, CLK=>clk, 
      R=>rst);
   ix10385 : aoi21 port map ( Y=>nx10384, A0=>label_5_output(0), A1=>nx35763, 
      B0=>nx36387);
   ix21584 : oai21 port map ( Y=>nx21583, A0=>nx29502, A1=>nx34765, B0=>
      nx29504);
   max_calc_reg_comparator_third_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx29502, D=>nx21583, CLK=>clk);
   ix29505 : nand03 port map ( Y=>nx29504, A0=>label_6_output(0), A1=>
      nx35453, A2=>nx34765);
   labelsregfile_label6_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_6_output(0), QB=>OPEN, D=>nx21033, CLK=>clk, R=>rst);
   lat_label_6_input_0 : latch port map ( Q=>label_6_input_0, D=>nx11718, 
      CLK=>nx34521);
   ix11719 : oai21 port map ( Y=>nx11718, A0=>nx29510, A1=>nx34419, B0=>
      nx29514);
   reg_label_6_input_state_machine_0 : dffr port map ( Q=>
      label_6_input_state_machine_0, QB=>nx29510, D=>nx21023, CLK=>clk, R=>
      rst);
   ix29515 : oai21 port map ( Y=>nx29514, A0=>nx35767, A1=>label_6_output(0), 
      B0=>nx11706);
   booth_booth_integrtaion_5_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_1, QB=>OPEN, D=>nx21003, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_2, QB=>nx29935, D=>nx20993, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_3, QB=>OPEN, D=>nx20983, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_4, QB=>nx29933, D=>nx20973, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_5, QB=>OPEN, D=>nx20963, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_6, QB=>nx29931, D=>nx20953, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_7, QB=>OPEN, D=>nx20943, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_8, QB=>nx29929, D=>nx20933, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_9, QB=>OPEN, D=>nx20923, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_10, QB=>nx29927, D=>nx20913, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_11, QB=>OPEN, D=>nx20903, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_12, QB=>nx29925, D=>nx20893, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_13, QB=>OPEN, D=>nx20883, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_14, QB=>nx29923, D=>nx20873, CLK=>clk, 
      R=>rst);
   ix29564 : aoi22 port map ( Y=>nx29563, A0=>mdr_data_out(15), A1=>nx34971, 
      B0=>nx11504, B1=>nx11510);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_reg_output_0, QB=>OPEN, 
      D=>nx20513, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_0, QB=>OPEN, D=>nx20499, CLK
      =>clk, S=>nx34483);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_reg_output_9, QB=>OPEN, 
      D=>nx20693, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_9, QB=>OPEN, D=>nx20683, CLK
      =>clk, R=>nx34483);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_8, QB=>OPEN, 
      D=>nx20673, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_8, QB=>OPEN, D=>nx20663, CLK
      =>clk, R=>nx34483);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_7, QB=>OPEN, 
      D=>nx20653, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_7, QB=>OPEN, D=>nx20643, CLK
      =>clk, R=>nx34483);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_6, QB=>OPEN, 
      D=>nx20633, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_6, QB=>OPEN, D=>nx20623, CLK
      =>clk, R=>nx34483);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_5, QB=>OPEN, 
      D=>nx20613, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_5, QB=>OPEN, D=>nx20603, CLK
      =>clk, R=>nx34483);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_4, QB=>OPEN, 
      D=>nx20593, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_4, QB=>OPEN, D=>nx20583, CLK
      =>clk, R=>nx34481);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_3, QB=>OPEN, 
      D=>nx20573, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_3, QB=>OPEN, D=>nx20563, CLK
      =>clk, R=>nx34481);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_2, QB=>OPEN, 
      D=>nx20553, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_2, QB=>OPEN, D=>nx20543, CLK
      =>clk, R=>nx34481);
   booth_booth_integrtaion_5_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_5_shift_Reg_output_1, QB=>OPEN, 
      D=>nx20533, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_5_shift_Reg_count_1, QB=>OPEN, D=>nx20523, CLK
      =>clk, R=>nx34481);
   ix20494 : nand02 port map ( Y=>nx20493, A0=>nx35827, A1=>nx34957);
   booth_booth_integrtaion_5_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx29610, D=>nx20493, CLK=>clk, S=>nx34481);
   ix11505 : nand02 port map ( Y=>nx11504, A0=>nx29631, A1=>nx29643);
   ix29632 : oai21 port map ( Y=>nx29631, A0=>nx34985, A1=>nx34979, B0=>
      mdr_data_out(96));
   ix20704 : oai21 port map ( Y=>nx20703, A0=>nx29636, A1=>nx35473, B0=>
      nx29638);
   booth_booth_integrtaion_5_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx29636, D=>nx20703, CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx29640, D=>nx21013, CLK=>clk, R=>rst);
   ix29648 : xnor2 port map ( Y=>nx29647, A0=>nx10974, A1=>nx13257);
   ix20844 : oai21 port map ( Y=>nx20843, A0=>nx29653, A1=>nx35473, B0=>
      nx29655);
   booth_booth_integrtaion_5_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_17, QB=>nx29653, D=>nx20843, 
      CLK=>clk, R=>rst);
   ix29656 : nand03 port map ( Y=>nx29655, A0=>nx35481, A1=>nx11482, A2=>
      nx36131);
   ix11483 : xnor2 port map ( Y=>nx11482, A0=>nx29658, A1=>nx13259);
   ix29659 : aoi22 port map ( Y=>nx29658, A0=>
      booth_booth_integrtaion_5_booth_output_17, A1=>nx10998, B0=>nx10974, 
      B1=>nx13257);
   ix10983 : nand02 port map ( Y=>nx10982, A0=>mdr_data_out(97), A1=>
      mdr_data_out(96));
   ix29663 : or02 port map ( Y=>nx29662, A0=>mdr_data_out(96), A1=>
      mdr_data_out(97));
   ix29669 : xnor2 port map ( Y=>nx29668, A0=>nx11026, A1=>nx13260);
   ix11027 : oai22 port map ( Y=>nx11026, A0=>nx29658, A1=>nx29671, B0=>
      nx29678, B1=>nx35485);
   ix29674 : aoi32 port map ( Y=>nx29673, A0=>nx11008, A1=>nx34985, A2=>
      nx29676, B0=>mdr_data_out(98), B1=>nx34979);
   ix11009 : oai21 port map ( Y=>nx11008, A0=>mdr_data_out(96), A1=>
      mdr_data_out(97), B0=>mdr_data_out(98));
   booth_booth_integrtaion_5_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_18, QB=>nx29678, D=>nx20833, 
      CLK=>clk, R=>rst);
   ix20824 : oai21 port map ( Y=>nx20823, A0=>nx29683, A1=>nx35473, B0=>
      nx29685);
   booth_booth_integrtaion_5_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_19, QB=>nx29683, D=>nx20823, 
      CLK=>clk, R=>rst);
   ix29686 : nand03 port map ( Y=>nx29685, A0=>nx35481, A1=>nx11458, A2=>
      nx36131);
   ix11459 : xnor2 port map ( Y=>nx11458, A0=>nx29688, A1=>nx13261);
   ix29689 : aoi22 port map ( Y=>nx29688, A0=>
      booth_booth_integrtaion_5_booth_output_19, A1=>nx11046, B0=>nx11026, 
      B1=>nx13260);
   ix29692 : nor02ii port map ( Y=>nx29691, A0=>nx11012, A1=>
      mdr_data_out(99));
   ix11013 : nor03_2x port map ( Y=>nx11012, A0=>mdr_data_out(98), A1=>
      mdr_data_out(96), A2=>mdr_data_out(97));
   ix11037 : nor04 port map ( Y=>nx11036, A0=>mdr_data_out(99), A1=>
      mdr_data_out(98), A2=>mdr_data_out(96), A3=>mdr_data_out(97));
   ix29706 : xnor2 port map ( Y=>nx29705, A0=>nx11074, A1=>nx13262);
   ix11075 : oai22 port map ( Y=>nx11074, A0=>nx29688, A1=>nx29708, B0=>
      nx29717, B1=>nx35487);
   ix29711 : aoi32 port map ( Y=>nx29710, A0=>nx11056, A1=>nx34985, A2=>
      nx29715, B0=>mdr_data_out(100), B1=>nx34979);
   ix11057 : nand02 port map ( Y=>nx11056, A0=>nx29713, A1=>
      mdr_data_out(100));
   booth_booth_integrtaion_5_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_20, QB=>nx29717, D=>nx20813, 
      CLK=>clk, R=>rst);
   ix20804 : oai21 port map ( Y=>nx20803, A0=>nx29722, A1=>nx35473, B0=>
      nx29724);
   booth_booth_integrtaion_5_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_21, QB=>nx29722, D=>nx20803, 
      CLK=>clk, R=>rst);
   ix29725 : nand03 port map ( Y=>nx29724, A0=>nx35481, A1=>nx11434, A2=>
      nx36131);
   ix11435 : xnor2 port map ( Y=>nx11434, A0=>nx29727, A1=>nx13263);
   ix29728 : aoi22 port map ( Y=>nx29727, A0=>
      booth_booth_integrtaion_5_booth_output_21, A1=>nx11094, B0=>nx11074, 
      B1=>nx13262);
   ix29731 : nor02ii port map ( Y=>nx29730, A0=>nx11060, A1=>
      mdr_data_out(101));
   ix11061 : nor02ii port map ( Y=>nx11060, A0=>mdr_data_out(100), A1=>
      nx11036);
   ix11085 : nor02ii port map ( Y=>nx11084, A0=>mdr_data_out(101), A1=>
      nx11060);
   ix29741 : xnor2 port map ( Y=>nx29740, A0=>nx11122, A1=>nx13264);
   ix11123 : oai22 port map ( Y=>nx11122, A0=>nx29727, A1=>nx29743, B0=>
      nx29752, B1=>nx35489);
   ix29746 : aoi32 port map ( Y=>nx29745, A0=>nx11104, A1=>nx34985, A2=>
      nx29750, B0=>mdr_data_out(102), B1=>nx34979);
   ix11105 : nand02 port map ( Y=>nx11104, A0=>nx29748, A1=>
      mdr_data_out(102));
   booth_booth_integrtaion_5_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_22, QB=>nx29752, D=>nx20793, 
      CLK=>clk, R=>rst);
   ix20784 : oai21 port map ( Y=>nx20783, A0=>nx29757, A1=>nx35473, B0=>
      nx29759);
   booth_booth_integrtaion_5_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_23, QB=>nx29757, D=>nx20783, 
      CLK=>clk, R=>rst);
   ix29760 : nand03 port map ( Y=>nx29759, A0=>nx35481, A1=>nx11410, A2=>
      nx35475);
   ix11411 : xnor2 port map ( Y=>nx11410, A0=>nx29762, A1=>nx13265);
   ix29763 : aoi22 port map ( Y=>nx29762, A0=>
      booth_booth_integrtaion_5_booth_output_23, A1=>nx11142, B0=>nx11122, 
      B1=>nx13264);
   ix29766 : nor02ii port map ( Y=>nx29765, A0=>nx11108, A1=>
      mdr_data_out(103));
   ix11109 : nor02ii port map ( Y=>nx11108, A0=>mdr_data_out(102), A1=>
      nx11084);
   ix11133 : nor02ii port map ( Y=>nx11132, A0=>mdr_data_out(103), A1=>
      nx11108);
   ix29776 : xnor2 port map ( Y=>nx29775, A0=>nx11170, A1=>nx13267);
   ix11171 : oai22 port map ( Y=>nx11170, A0=>nx29762, A1=>nx29778, B0=>
      nx29787, B1=>nx35491);
   ix29781 : aoi32 port map ( Y=>nx29780, A0=>nx11152, A1=>nx34985, A2=>
      nx29785, B0=>mdr_data_out(104), B1=>nx34979);
   ix11153 : nand02 port map ( Y=>nx11152, A0=>nx29783, A1=>
      mdr_data_out(104));
   booth_booth_integrtaion_5_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_24, QB=>nx29787, D=>nx20773, 
      CLK=>clk, R=>rst);
   ix20764 : oai21 port map ( Y=>nx20763, A0=>nx29792, A1=>nx35475, B0=>
      nx29794);
   booth_booth_integrtaion_5_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_25, QB=>nx29792, D=>nx20763, 
      CLK=>clk, R=>rst);
   ix29795 : nand03 port map ( Y=>nx29794, A0=>nx35481, A1=>nx11386, A2=>
      nx35475);
   ix11387 : xnor2 port map ( Y=>nx11386, A0=>nx29797, A1=>nx13269);
   ix29798 : aoi22 port map ( Y=>nx29797, A0=>
      booth_booth_integrtaion_5_booth_output_25, A1=>nx11190, B0=>nx11170, 
      B1=>nx13267);
   ix29801 : nor02ii port map ( Y=>nx29800, A0=>nx11156, A1=>
      mdr_data_out(105));
   ix11157 : nor02ii port map ( Y=>nx11156, A0=>mdr_data_out(104), A1=>
      nx11132);
   ix11181 : nor02ii port map ( Y=>nx11180, A0=>mdr_data_out(105), A1=>
      nx11156);
   ix29811 : xnor2 port map ( Y=>nx29810, A0=>nx11218, A1=>nx13271);
   ix11219 : oai22 port map ( Y=>nx11218, A0=>nx29797, A1=>nx29813, B0=>
      nx29822, B1=>nx35493);
   ix29816 : aoi32 port map ( Y=>nx29815, A0=>nx11200, A1=>nx34985, A2=>
      nx29820, B0=>mdr_data_out(106), B1=>nx34979);
   ix11201 : nand02 port map ( Y=>nx11200, A0=>nx29818, A1=>
      mdr_data_out(106));
   booth_booth_integrtaion_5_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_26, QB=>nx29822, D=>nx20753, 
      CLK=>clk, R=>rst);
   ix20744 : oai21 port map ( Y=>nx20743, A0=>nx29827, A1=>nx35475, B0=>
      nx29829);
   booth_booth_integrtaion_5_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_27, QB=>nx29827, D=>nx20743, 
      CLK=>clk, R=>rst);
   ix29830 : nand03 port map ( Y=>nx29829, A0=>nx35481, A1=>nx11362, A2=>
      nx35475);
   ix11363 : xnor2 port map ( Y=>nx11362, A0=>nx29832, A1=>nx13272);
   ix29833 : aoi22 port map ( Y=>nx29832, A0=>
      booth_booth_integrtaion_5_booth_output_27, A1=>nx11238, B0=>nx11218, 
      B1=>nx13271);
   ix29836 : nor02ii port map ( Y=>nx29835, A0=>nx11204, A1=>
      mdr_data_out(107));
   ix11205 : nor02ii port map ( Y=>nx11204, A0=>mdr_data_out(106), A1=>
      nx11180);
   ix11229 : nor02ii port map ( Y=>nx11228, A0=>mdr_data_out(107), A1=>
      nx11204);
   ix29846 : xnor2 port map ( Y=>nx29845, A0=>nx11266, A1=>nx13273);
   ix11267 : oai22 port map ( Y=>nx11266, A0=>nx29832, A1=>nx29848, B0=>
      nx29857, B1=>nx35495);
   ix29851 : aoi32 port map ( Y=>nx29850, A0=>nx11248, A1=>nx34985, A2=>
      nx29855, B0=>mdr_data_out(108), B1=>nx34979);
   ix11249 : nand02 port map ( Y=>nx11248, A0=>nx29853, A1=>
      mdr_data_out(108));
   booth_booth_integrtaion_5_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_28, QB=>nx29857, D=>nx20733, 
      CLK=>clk, R=>rst);
   ix20724 : oai21 port map ( Y=>nx20723, A0=>nx29862, A1=>nx35475, B0=>
      nx29864);
   booth_booth_integrtaion_5_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_29, QB=>nx29862, D=>nx20723, 
      CLK=>clk, R=>rst);
   ix29865 : nand03 port map ( Y=>nx29864, A0=>nx36139, A1=>nx11338, A2=>
      nx35475);
   ix11339 : xnor2 port map ( Y=>nx11338, A0=>nx29867, A1=>nx13274);
   ix29868 : aoi22 port map ( Y=>nx29867, A0=>
      booth_booth_integrtaion_5_booth_output_29, A1=>nx11286, B0=>nx11266, 
      B1=>nx13273);
   ix29871 : nor02ii port map ( Y=>nx29870, A0=>nx11252, A1=>
      mdr_data_out(109));
   ix11253 : nor02ii port map ( Y=>nx11252, A0=>mdr_data_out(108), A1=>
      nx11228);
   ix11277 : nor02ii port map ( Y=>nx11276, A0=>mdr_data_out(109), A1=>
      nx11252);
   ix29881 : xnor2 port map ( Y=>nx29880, A0=>nx11314, A1=>nx11324);
   ix11315 : oai22 port map ( Y=>nx11314, A0=>nx29867, A1=>nx29883, B0=>
      nx29892, B1=>nx35497);
   ix29886 : aoi32 port map ( Y=>nx29885, A0=>nx11296, A1=>nx34987, A2=>
      nx29890, B0=>mdr_data_out(110), B1=>nx34981);
   ix11297 : nand02 port map ( Y=>nx11296, A0=>nx29888, A1=>
      mdr_data_out(110));
   booth_booth_integrtaion_5_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_31, QB=>nx29892, D=>nx20713, 
      CLK=>clk, R=>rst);
   ix29896 : aoi22 port map ( Y=>nx29895, A0=>mdr_data_out(111), A1=>nx34981, 
      B0=>nx34987, B1=>nx11316);
   ix11317 : xnor2 port map ( Y=>nx11316, A0=>mdr_data_out(111), A1=>nx11300
   );
   ix11301 : nor02ii port map ( Y=>nx11300, A0=>mdr_data_out(110), A1=>
      nx11276);
   ix29900 : aoi32 port map ( Y=>nx29899, A0=>nx11272, A1=>nx34987, A2=>
      nx29888, B0=>mdr_data_out(109), B1=>nx34981);
   ix29903 : aoi32 port map ( Y=>nx29902, A0=>nx11224, A1=>nx34987, A2=>
      nx29853, B0=>mdr_data_out(107), B1=>nx34981);
   ix29906 : aoi32 port map ( Y=>nx29905, A0=>nx11176, A1=>nx34987, A2=>
      nx29818, B0=>mdr_data_out(105), B1=>nx34981);
   ix29909 : aoi32 port map ( Y=>nx29908, A0=>nx11128, A1=>nx34987, A2=>
      nx29783, B0=>mdr_data_out(103), B1=>nx34981);
   ix29912 : aoi32 port map ( Y=>nx29911, A0=>nx11080, A1=>nx34987, A2=>
      nx29748, B0=>mdr_data_out(101), B1=>nx34981);
   ix29915 : aoi32 port map ( Y=>nx29914, A0=>nx11032, A1=>nx10968, A2=>
      nx29713, B0=>mdr_data_out(99), B1=>nx34983);
   ix29918 : aoi32 port map ( Y=>nx29917, A0=>nx10982, A1=>nx10968, A2=>
      nx29662, B0=>mdr_data_out(97), B1=>nx34983);
   booth_booth_integrtaion_5_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_5_booth_output_16, QB=>nx29643, D=>nx20853, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_5_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_5_15, QB=>nx29921, D=>nx20863, CLK=>clk, 
      R=>rst);
   ix11707 : aoi21 port map ( Y=>nx11706, A0=>label_6_output(0), A1=>nx35767, 
      B0=>nx36387);
   ix12691 : xnor2 port map ( Y=>nx12690, A0=>nx29940, A1=>nx12688);
   ix29941 : aoi22 port map ( Y=>nx29940, A0=>nx29942, A1=>
      max_calc_comparator_third_inp1_14, B0=>nx12176, B1=>nx12594);
   max_calc_reg_comparator_third_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx29942, D=>nx21313, CLK=>clk);
   ix21314 : oai21 port map ( Y=>nx21313, A0=>nx29942, A1=>nx34765, B0=>
      nx29945);
   labelsregfile_label6_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_6_output(14), QB=>nx30129, D=>nx21303, CLK=>clk, R=>rst);
   lat_label_6_input_14 : latch port map ( Q=>label_6_input_14, D=>nx12154, 
      CLK=>nx34525);
   reg_label_6_input_state_machine_14 : dffr port map ( Q=>
      label_6_input_state_machine_14, QB=>OPEN, D=>nx20483, CLK=>clk, R=>rst
   );
   ix12151 : xor2 port map ( Y=>nx12150, A0=>nx29955, A1=>nx30127);
   ix29956 : aoi22 port map ( Y=>nx29955, A0=>label_6_output(13), A1=>
      booth_booth_integration_output_5_13, B0=>nx12114, B1=>nx13293);
   labelsregfile_label6_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_6_output(13), QB=>OPEN, D=>nx21293, CLK=>clk, R=>rst);
   lat_label_6_input_13 : latch port map ( Q=>label_6_input_13, D=>nx12128, 
      CLK=>nx34525);
   reg_label_6_input_state_machine_13 : dffr port map ( Q=>
      label_6_input_state_machine_13, QB=>OPEN, D=>nx21283, CLK=>clk, R=>rst
   );
   ix12125 : xnor2 port map ( Y=>nx12124, A0=>nx12114, A1=>nx30123);
   ix12115 : oai22 port map ( Y=>nx12114, A0=>nx29966, A1=>nx30112, B0=>
      nx30122, B1=>nx29925);
   ix29967 : aoi22 port map ( Y=>nx29966, A0=>label_6_output(11), A1=>
      booth_booth_integration_output_5_11, B0=>nx12050, B1=>nx13289);
   labelsregfile_label6_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_6_output(11), QB=>OPEN, D=>nx21253, CLK=>clk, R=>rst);
   lat_label_6_input_11 : latch port map ( Q=>label_6_input_11, D=>nx12064, 
      CLK=>nx34523);
   reg_label_6_input_state_machine_11 : dffr port map ( Q=>
      label_6_input_state_machine_11, QB=>OPEN, D=>nx21243, CLK=>clk, R=>rst
   );
   ix12061 : xnor2 port map ( Y=>nx12060, A0=>nx12050, A1=>nx30108);
   ix12051 : oai22 port map ( Y=>nx12050, A0=>nx29977, A1=>nx30097, B0=>
      nx30107, B1=>nx29927);
   ix29978 : aoi22 port map ( Y=>nx29977, A0=>label_6_output(9), A1=>
      booth_booth_integration_output_5_9, B0=>nx11986, B1=>nx13287);
   labelsregfile_label6_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_6_output(9), QB=>OPEN, D=>nx21213, CLK=>clk, R=>rst);
   lat_label_6_input_9 : latch port map ( Q=>label_6_input_9, D=>nx12000, 
      CLK=>nx34523);
   reg_label_6_input_state_machine_9 : dffr port map ( Q=>
      label_6_input_state_machine_9, QB=>OPEN, D=>nx21203, CLK=>clk, R=>rst
   );
   ix11997 : xnor2 port map ( Y=>nx11996, A0=>nx11986, A1=>nx30093);
   ix11987 : oai22 port map ( Y=>nx11986, A0=>nx29988, A1=>nx30082, B0=>
      nx30092, B1=>nx29929);
   ix29989 : aoi22 port map ( Y=>nx29988, A0=>label_6_output(7), A1=>
      booth_booth_integration_output_5_7, B0=>nx11922, B1=>nx13285);
   labelsregfile_label6_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_6_output(7), QB=>OPEN, D=>nx21173, CLK=>clk, R=>rst);
   lat_label_6_input_7 : latch port map ( Q=>label_6_input_7, D=>nx11936, 
      CLK=>nx34523);
   reg_label_6_input_state_machine_7 : dffr port map ( Q=>
      label_6_input_state_machine_7, QB=>OPEN, D=>nx21163, CLK=>clk, R=>rst
   );
   ix11933 : xnor2 port map ( Y=>nx11932, A0=>nx11922, A1=>nx30078);
   ix11923 : oai22 port map ( Y=>nx11922, A0=>nx29999, A1=>nx30067, B0=>
      nx30077, B1=>nx29931);
   ix30000 : aoi22 port map ( Y=>nx29999, A0=>label_6_output(5), A1=>
      booth_booth_integration_output_5_5, B0=>nx11858, B1=>nx13283);
   labelsregfile_label6_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_6_output(5), QB=>OPEN, D=>nx21133, CLK=>clk, R=>rst);
   lat_label_6_input_5 : latch port map ( Q=>label_6_input_5, D=>nx11872, 
      CLK=>nx34521);
   reg_label_6_input_state_machine_5 : dffr port map ( Q=>
      label_6_input_state_machine_5, QB=>OPEN, D=>nx21123, CLK=>clk, R=>rst
   );
   ix11869 : xnor2 port map ( Y=>nx11868, A0=>nx11858, A1=>nx30063);
   ix11859 : oai22 port map ( Y=>nx11858, A0=>nx30010, A1=>nx30052, B0=>
      nx30062, B1=>nx29933);
   ix30011 : aoi22 port map ( Y=>nx30010, A0=>label_6_output(3), A1=>
      booth_booth_integration_output_5_3, B0=>nx11794, B1=>nx13279);
   labelsregfile_label6_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_6_output(3), QB=>OPEN, D=>nx21093, CLK=>clk, R=>rst);
   lat_label_6_input_3 : latch port map ( Q=>label_6_input_3, D=>nx11808, 
      CLK=>nx34521);
   reg_label_6_input_state_machine_3 : dffr port map ( Q=>
      label_6_input_state_machine_3, QB=>OPEN, D=>nx21083, CLK=>clk, R=>rst
   );
   ix11805 : xnor2 port map ( Y=>nx11804, A0=>nx11794, A1=>nx30048);
   ix11795 : oai22 port map ( Y=>nx11794, A0=>nx30021, A1=>nx30037, B0=>
      nx30047, B1=>nx29935);
   ix30022 : aoi32 port map ( Y=>nx30021, A0=>label_6_output(0), A1=>nx35767, 
      A2=>nx13276, B0=>label_6_output(1), B1=>
      booth_booth_integration_output_5_1);
   labelsregfile_label6_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_6_output(1), QB=>OPEN, D=>nx21053, CLK=>clk, R=>rst);
   lat_label_6_input_1 : latch port map ( Q=>label_6_input_1, D=>nx11744, 
      CLK=>nx34521);
   reg_label_6_input_state_machine_1 : dffr port map ( Q=>
      label_6_input_state_machine_1, QB=>OPEN, D=>nx21043, CLK=>clk, R=>rst
   );
   ix11741 : xor2 port map ( Y=>nx11740, A0=>nx30032, A1=>nx30034);
   ix30033 : nand02 port map ( Y=>nx30032, A0=>label_6_output(0), A1=>
      nx35767);
   ix30035 : xnor2 port map ( Y=>nx30034, A0=>
      booth_booth_integration_output_5_1, A1=>label_6_output(1));
   labelsregfile_label6_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_6_output(2), QB=>nx30047, D=>nx21073, CLK=>clk, R=>rst);
   lat_label_6_input_2 : latch port map ( Q=>label_6_input_2, D=>nx11776, 
      CLK=>nx34521);
   reg_label_6_input_state_machine_2 : dffr port map ( Q=>
      label_6_input_state_machine_2, QB=>OPEN, D=>nx21063, CLK=>clk, R=>rst
   );
   ix11773 : xor2 port map ( Y=>nx11772, A0=>nx30021, A1=>nx30037);
   ix30049 : xnor2 port map ( Y=>nx30048, A0=>
      booth_booth_integration_output_5_3, A1=>label_6_output(3));
   labelsregfile_label6_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_6_output(4), QB=>nx30062, D=>nx21113, CLK=>clk, R=>rst);
   lat_label_6_input_4 : latch port map ( Q=>label_6_input_4, D=>nx11840, 
      CLK=>nx34521);
   reg_label_6_input_state_machine_4 : dffr port map ( Q=>
      label_6_input_state_machine_4, QB=>OPEN, D=>nx21103, CLK=>clk, R=>rst
   );
   ix11837 : xor2 port map ( Y=>nx11836, A0=>nx30010, A1=>nx30052);
   ix30064 : xnor2 port map ( Y=>nx30063, A0=>
      booth_booth_integration_output_5_5, A1=>label_6_output(5));
   labelsregfile_label6_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_6_output(6), QB=>nx30077, D=>nx21153, CLK=>clk, R=>rst);
   lat_label_6_input_6 : latch port map ( Q=>label_6_input_6, D=>nx11904, 
      CLK=>nx34523);
   reg_label_6_input_state_machine_6 : dffr port map ( Q=>
      label_6_input_state_machine_6, QB=>OPEN, D=>nx21143, CLK=>clk, R=>rst
   );
   ix11901 : xor2 port map ( Y=>nx11900, A0=>nx29999, A1=>nx30067);
   ix30079 : xnor2 port map ( Y=>nx30078, A0=>
      booth_booth_integration_output_5_7, A1=>label_6_output(7));
   labelsregfile_label6_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_6_output(8), QB=>nx30092, D=>nx21193, CLK=>clk, R=>rst);
   lat_label_6_input_8 : latch port map ( Q=>label_6_input_8, D=>nx11968, 
      CLK=>nx34523);
   reg_label_6_input_state_machine_8 : dffr port map ( Q=>
      label_6_input_state_machine_8, QB=>OPEN, D=>nx21183, CLK=>clk, R=>rst
   );
   ix11965 : xor2 port map ( Y=>nx11964, A0=>nx29988, A1=>nx30082);
   ix30094 : xnor2 port map ( Y=>nx30093, A0=>
      booth_booth_integration_output_5_9, A1=>label_6_output(9));
   labelsregfile_label6_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_6_output(10), QB=>nx30107, D=>nx21233, CLK=>clk, R=>rst);
   lat_label_6_input_10 : latch port map ( Q=>label_6_input_10, D=>nx12032, 
      CLK=>nx34523);
   reg_label_6_input_state_machine_10 : dffr port map ( Q=>
      label_6_input_state_machine_10, QB=>OPEN, D=>nx21223, CLK=>clk, R=>rst
   );
   ix12029 : xor2 port map ( Y=>nx12028, A0=>nx29977, A1=>nx30097);
   ix30109 : xnor2 port map ( Y=>nx30108, A0=>
      booth_booth_integration_output_5_11, A1=>label_6_output(11));
   labelsregfile_label6_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_6_output(12), QB=>nx30122, D=>nx21273, CLK=>clk, R=>rst);
   lat_label_6_input_12 : latch port map ( Q=>label_6_input_12, D=>nx12096, 
      CLK=>nx34523);
   reg_label_6_input_state_machine_12 : dffr port map ( Q=>
      label_6_input_state_machine_12, QB=>OPEN, D=>nx21263, CLK=>clk, R=>rst
   );
   ix12093 : xor2 port map ( Y=>nx12092, A0=>nx29966, A1=>nx30112);
   ix30124 : xnor2 port map ( Y=>nx30123, A0=>
      booth_booth_integration_output_5_13, A1=>label_6_output(13));
   ix20474 : oai21 port map ( Y=>nx20473, A0=>nx30132, A1=>nx34767, B0=>
      nx30134);
   max_calc_reg_comparator_third_inp1_14 : dff port map ( Q=>
      max_calc_comparator_third_inp1_14, QB=>nx30132, D=>nx20473, CLK=>clk);
   labelsregfile_label5_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_5_output(14), QB=>nx30318, D=>nx20463, CLK=>clk, R=>rst);
   lat_label_5_input_14 : latch port map ( Q=>label_5_input_14, D=>nx10832, 
      CLK=>nx34529);
   reg_label_5_input_state_machine_14 : dffr port map ( Q=>
      label_5_input_state_machine_14, QB=>OPEN, D=>nx19643, CLK=>clk, R=>rst
   );
   ix10829 : xor2 port map ( Y=>nx10828, A0=>nx30144, A1=>nx30316);
   ix30145 : aoi22 port map ( Y=>nx30144, A0=>label_5_output(13), A1=>
      booth_booth_integration_output_4_13, B0=>nx10792, B1=>nx13253);
   labelsregfile_label5_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_5_output(13), QB=>OPEN, D=>nx20453, CLK=>clk, R=>rst);
   lat_label_5_input_13 : latch port map ( Q=>label_5_input_13, D=>nx10806, 
      CLK=>nx34529);
   reg_label_5_input_state_machine_13 : dffr port map ( Q=>
      label_5_input_state_machine_13, QB=>OPEN, D=>nx20443, CLK=>clk, R=>rst
   );
   ix10803 : xnor2 port map ( Y=>nx10802, A0=>nx10792, A1=>nx30312);
   ix10793 : oai22 port map ( Y=>nx10792, A0=>nx30155, A1=>nx30301, B0=>
      nx30311, B1=>nx29484);
   ix30156 : aoi22 port map ( Y=>nx30155, A0=>label_5_output(11), A1=>
      booth_booth_integration_output_4_11, B0=>nx10728, B1=>nx13251);
   labelsregfile_label5_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_5_output(11), QB=>OPEN, D=>nx20413, CLK=>clk, R=>rst);
   lat_label_5_input_11 : latch port map ( Q=>label_5_input_11, D=>nx10742, 
      CLK=>nx34527);
   reg_label_5_input_state_machine_11 : dffr port map ( Q=>
      label_5_input_state_machine_11, QB=>OPEN, D=>nx20403, CLK=>clk, R=>rst
   );
   ix10739 : xnor2 port map ( Y=>nx10738, A0=>nx10728, A1=>nx30297);
   ix10729 : oai22 port map ( Y=>nx10728, A0=>nx30166, A1=>nx30286, B0=>
      nx30296, B1=>nx29486);
   ix30167 : aoi22 port map ( Y=>nx30166, A0=>label_5_output(9), A1=>
      booth_booth_integration_output_4_9, B0=>nx10664, B1=>nx13249);
   labelsregfile_label5_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_5_output(9), QB=>OPEN, D=>nx20373, CLK=>clk, R=>rst);
   lat_label_5_input_9 : latch port map ( Q=>label_5_input_9, D=>nx10678, 
      CLK=>nx34527);
   reg_label_5_input_state_machine_9 : dffr port map ( Q=>
      label_5_input_state_machine_9, QB=>OPEN, D=>nx20363, CLK=>clk, R=>rst
   );
   ix10675 : xnor2 port map ( Y=>nx10674, A0=>nx10664, A1=>nx30282);
   ix10665 : oai22 port map ( Y=>nx10664, A0=>nx30177, A1=>nx30271, B0=>
      nx30281, B1=>nx29488);
   ix30178 : aoi22 port map ( Y=>nx30177, A0=>label_5_output(7), A1=>
      booth_booth_integration_output_4_7, B0=>nx10600, B1=>nx13247);
   labelsregfile_label5_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_5_output(7), QB=>OPEN, D=>nx20333, CLK=>clk, R=>rst);
   lat_label_5_input_7 : latch port map ( Q=>label_5_input_7, D=>nx10614, 
      CLK=>nx34527);
   reg_label_5_input_state_machine_7 : dffr port map ( Q=>
      label_5_input_state_machine_7, QB=>OPEN, D=>nx20323, CLK=>clk, R=>rst
   );
   ix10611 : xnor2 port map ( Y=>nx10610, A0=>nx10600, A1=>nx30267);
   ix10601 : oai22 port map ( Y=>nx10600, A0=>nx30188, A1=>nx30256, B0=>
      nx30266, B1=>nx29490);
   ix30189 : aoi22 port map ( Y=>nx30188, A0=>label_5_output(5), A1=>
      booth_booth_integration_output_4_5, B0=>nx10536, B1=>nx13243);
   labelsregfile_label5_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_5_output(5), QB=>OPEN, D=>nx20293, CLK=>clk, R=>rst);
   lat_label_5_input_5 : latch port map ( Q=>label_5_input_5, D=>nx10550, 
      CLK=>nx34525);
   reg_label_5_input_state_machine_5 : dffr port map ( Q=>
      label_5_input_state_machine_5, QB=>OPEN, D=>nx20283, CLK=>clk, R=>rst
   );
   ix10547 : xnor2 port map ( Y=>nx10546, A0=>nx10536, A1=>nx30252);
   ix10537 : oai22 port map ( Y=>nx10536, A0=>nx30199, A1=>nx30241, B0=>
      nx30251, B1=>nx29492);
   ix30200 : aoi22 port map ( Y=>nx30199, A0=>label_5_output(3), A1=>
      booth_booth_integration_output_4_3, B0=>nx10472, B1=>nx13240);
   labelsregfile_label5_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_5_output(3), QB=>OPEN, D=>nx20253, CLK=>clk, R=>rst);
   lat_label_5_input_3 : latch port map ( Q=>label_5_input_3, D=>nx10486, 
      CLK=>nx34525);
   reg_label_5_input_state_machine_3 : dffr port map ( Q=>
      label_5_input_state_machine_3, QB=>OPEN, D=>nx20243, CLK=>clk, R=>rst
   );
   ix10483 : xnor2 port map ( Y=>nx10482, A0=>nx10472, A1=>nx30237);
   ix10473 : oai22 port map ( Y=>nx10472, A0=>nx30210, A1=>nx30226, B0=>
      nx30236, B1=>nx29494);
   ix30211 : aoi32 port map ( Y=>nx30210, A0=>label_5_output(0), A1=>nx35763, 
      A2=>nx13238, B0=>label_5_output(1), B1=>
      booth_booth_integration_output_4_1);
   labelsregfile_label5_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_5_output(1), QB=>OPEN, D=>nx20213, CLK=>clk, R=>rst);
   lat_label_5_input_1 : latch port map ( Q=>label_5_input_1, D=>nx10422, 
      CLK=>nx34525);
   reg_label_5_input_state_machine_1 : dffr port map ( Q=>
      label_5_input_state_machine_1, QB=>OPEN, D=>nx20203, CLK=>clk, R=>rst
   );
   ix10419 : xor2 port map ( Y=>nx10418, A0=>nx30221, A1=>nx30223);
   ix30222 : nand02 port map ( Y=>nx30221, A0=>label_5_output(0), A1=>
      nx35763);
   ix30224 : xnor2 port map ( Y=>nx30223, A0=>
      booth_booth_integration_output_4_1, A1=>label_5_output(1));
   labelsregfile_label5_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_5_output(2), QB=>nx30236, D=>nx20233, CLK=>clk, R=>rst);
   lat_label_5_input_2 : latch port map ( Q=>label_5_input_2, D=>nx10454, 
      CLK=>nx34525);
   reg_label_5_input_state_machine_2 : dffr port map ( Q=>
      label_5_input_state_machine_2, QB=>OPEN, D=>nx20223, CLK=>clk, R=>rst
   );
   ix10451 : xor2 port map ( Y=>nx10450, A0=>nx30210, A1=>nx30226);
   ix30238 : xnor2 port map ( Y=>nx30237, A0=>
      booth_booth_integration_output_4_3, A1=>label_5_output(3));
   labelsregfile_label5_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_5_output(4), QB=>nx30251, D=>nx20273, CLK=>clk, R=>rst);
   lat_label_5_input_4 : latch port map ( Q=>label_5_input_4, D=>nx10518, 
      CLK=>nx34525);
   reg_label_5_input_state_machine_4 : dffr port map ( Q=>
      label_5_input_state_machine_4, QB=>OPEN, D=>nx20263, CLK=>clk, R=>rst
   );
   ix10515 : xor2 port map ( Y=>nx10514, A0=>nx30199, A1=>nx30241);
   ix30253 : xnor2 port map ( Y=>nx30252, A0=>
      booth_booth_integration_output_4_5, A1=>label_5_output(5));
   labelsregfile_label5_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_5_output(6), QB=>nx30266, D=>nx20313, CLK=>clk, R=>rst);
   lat_label_5_input_6 : latch port map ( Q=>label_5_input_6, D=>nx10582, 
      CLK=>nx34527);
   reg_label_5_input_state_machine_6 : dffr port map ( Q=>
      label_5_input_state_machine_6, QB=>OPEN, D=>nx20303, CLK=>clk, R=>rst
   );
   ix10579 : xor2 port map ( Y=>nx10578, A0=>nx30188, A1=>nx30256);
   ix30268 : xnor2 port map ( Y=>nx30267, A0=>
      booth_booth_integration_output_4_7, A1=>label_5_output(7));
   labelsregfile_label5_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_5_output(8), QB=>nx30281, D=>nx20353, CLK=>clk, R=>rst);
   lat_label_5_input_8 : latch port map ( Q=>label_5_input_8, D=>nx10646, 
      CLK=>nx34527);
   reg_label_5_input_state_machine_8 : dffr port map ( Q=>
      label_5_input_state_machine_8, QB=>OPEN, D=>nx20343, CLK=>clk, R=>rst
   );
   ix10643 : xor2 port map ( Y=>nx10642, A0=>nx30177, A1=>nx30271);
   ix30283 : xnor2 port map ( Y=>nx30282, A0=>
      booth_booth_integration_output_4_9, A1=>label_5_output(9));
   labelsregfile_label5_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_5_output(10), QB=>nx30296, D=>nx20393, CLK=>clk, R=>rst);
   lat_label_5_input_10 : latch port map ( Q=>label_5_input_10, D=>nx10710, 
      CLK=>nx34527);
   reg_label_5_input_state_machine_10 : dffr port map ( Q=>
      label_5_input_state_machine_10, QB=>OPEN, D=>nx20383, CLK=>clk, R=>rst
   );
   ix10707 : xor2 port map ( Y=>nx10706, A0=>nx30166, A1=>nx30286);
   ix30298 : xnor2 port map ( Y=>nx30297, A0=>
      booth_booth_integration_output_4_11, A1=>label_5_output(11));
   labelsregfile_label5_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_5_output(12), QB=>nx30311, D=>nx20433, CLK=>clk, R=>rst);
   lat_label_5_input_12 : latch port map ( Q=>label_5_input_12, D=>nx10774, 
      CLK=>nx34527);
   reg_label_5_input_state_machine_12 : dffr port map ( Q=>
      label_5_input_state_machine_12, QB=>OPEN, D=>nx20423, CLK=>clk, R=>rst
   );
   ix10771 : xor2 port map ( Y=>nx10770, A0=>nx30155, A1=>nx30301);
   ix30313 : xnor2 port map ( Y=>nx30312, A0=>
      booth_booth_integration_output_4_13, A1=>label_5_output(13));
   ix12595 : oai22 port map ( Y=>nx12594, A0=>nx30321, A1=>nx30334, B0=>
      max_calc_comparator_third_inp2_13, B1=>nx30329);
   ix21324 : oai21 port map ( Y=>nx21323, A0=>nx30325, A1=>nx34767, B0=>
      nx30327);
   max_calc_reg_comparator_third_inp2_13 : dff port map ( Q=>
      max_calc_comparator_third_inp2_13, QB=>nx30325, D=>nx21323, CLK=>clk);
   ix30328 : nand03 port map ( Y=>nx30327, A0=>label_6_output(13), A1=>
      nx35453, A2=>nx34767);
   max_calc_reg_comparator_third_inp1_13 : dff port map ( Q=>
      max_calc_comparator_third_inp1_13, QB=>nx30329, D=>nx21333, CLK=>clk);
   ix21334 : oai21 port map ( Y=>nx21333, A0=>nx30329, A1=>nx34767, B0=>
      nx30332);
   ix30333 : nand03 port map ( Y=>nx30332, A0=>label_5_output(13), A1=>
      nx35453, A2=>nx34767);
   ix30335 : aoi22 port map ( Y=>nx30334, A0=>nx30336, A1=>
      max_calc_comparator_third_inp1_12, B0=>nx12220, B1=>nx12578);
   max_calc_reg_comparator_third_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx30336, D=>nx21343, CLK=>clk);
   ix21344 : oai21 port map ( Y=>nx21343, A0=>nx30336, A1=>nx34769, B0=>
      nx30339);
   ix21354 : oai21 port map ( Y=>nx21353, A0=>nx30343, A1=>nx34769, B0=>
      nx30345);
   max_calc_reg_comparator_third_inp1_12 : dff port map ( Q=>
      max_calc_comparator_third_inp1_12, QB=>nx30343, D=>nx21353, CLK=>clk);
   ix12579 : oai22 port map ( Y=>nx12578, A0=>nx30349, A1=>nx30362, B0=>
      max_calc_comparator_third_inp2_11, B1=>nx30357);
   ix21364 : oai21 port map ( Y=>nx21363, A0=>nx30353, A1=>nx34769, B0=>
      nx30355);
   max_calc_reg_comparator_third_inp2_11 : dff port map ( Q=>
      max_calc_comparator_third_inp2_11, QB=>nx30353, D=>nx21363, CLK=>clk);
   ix30356 : nand03 port map ( Y=>nx30355, A0=>label_6_output(11), A1=>
      nx35455, A2=>nx34769);
   max_calc_reg_comparator_third_inp1_11 : dff port map ( Q=>
      max_calc_comparator_third_inp1_11, QB=>nx30357, D=>nx21373, CLK=>clk);
   ix21374 : oai21 port map ( Y=>nx21373, A0=>nx30357, A1=>nx34769, B0=>
      nx30360);
   ix30361 : nand03 port map ( Y=>nx30360, A0=>label_5_output(11), A1=>
      nx35455, A2=>nx34771);
   ix30363 : aoi22 port map ( Y=>nx30362, A0=>nx30364, A1=>
      max_calc_comparator_third_inp1_10, B0=>nx12264, B1=>nx12562);
   max_calc_reg_comparator_third_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx30364, D=>nx21383, CLK=>clk);
   ix21384 : oai21 port map ( Y=>nx21383, A0=>nx30364, A1=>nx34771, B0=>
      nx30367);
   ix21394 : oai21 port map ( Y=>nx21393, A0=>nx30371, A1=>nx34771, B0=>
      nx30373);
   max_calc_reg_comparator_third_inp1_10 : dff port map ( Q=>
      max_calc_comparator_third_inp1_10, QB=>nx30371, D=>nx21393, CLK=>clk);
   ix12563 : oai22 port map ( Y=>nx12562, A0=>nx30377, A1=>nx30390, B0=>
      max_calc_comparator_third_inp2_9, B1=>nx30385);
   ix21404 : oai21 port map ( Y=>nx21403, A0=>nx30381, A1=>nx34771, B0=>
      nx30383);
   max_calc_reg_comparator_third_inp2_9 : dff port map ( Q=>
      max_calc_comparator_third_inp2_9, QB=>nx30381, D=>nx21403, CLK=>clk);
   ix30384 : nand03 port map ( Y=>nx30383, A0=>label_6_output(9), A1=>
      nx35455, A2=>nx34771);
   max_calc_reg_comparator_third_inp1_9 : dff port map ( Q=>
      max_calc_comparator_third_inp1_9, QB=>nx30385, D=>nx21413, CLK=>clk);
   ix21414 : oai21 port map ( Y=>nx21413, A0=>nx30385, A1=>nx34773, B0=>
      nx30388);
   ix30389 : nand03 port map ( Y=>nx30388, A0=>label_5_output(9), A1=>
      nx35455, A2=>nx34773);
   ix30391 : aoi22 port map ( Y=>nx30390, A0=>nx30392, A1=>
      max_calc_comparator_third_inp1_8, B0=>nx12308, B1=>nx12546);
   max_calc_reg_comparator_third_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx30392, D=>nx21423, CLK=>clk);
   ix21424 : oai21 port map ( Y=>nx21423, A0=>nx30392, A1=>nx34773, B0=>
      nx30395);
   ix21434 : oai21 port map ( Y=>nx21433, A0=>nx30399, A1=>nx34773, B0=>
      nx30401);
   max_calc_reg_comparator_third_inp1_8 : dff port map ( Q=>
      max_calc_comparator_third_inp1_8, QB=>nx30399, D=>nx21433, CLK=>clk);
   ix12547 : oai22 port map ( Y=>nx12546, A0=>nx30405, A1=>nx30418, B0=>
      max_calc_comparator_third_inp2_7, B1=>nx30413);
   ix21444 : oai21 port map ( Y=>nx21443, A0=>nx30409, A1=>nx34773, B0=>
      nx30411);
   max_calc_reg_comparator_third_inp2_7 : dff port map ( Q=>
      max_calc_comparator_third_inp2_7, QB=>nx30409, D=>nx21443, CLK=>clk);
   ix30412 : nand03 port map ( Y=>nx30411, A0=>label_6_output(7), A1=>
      nx35457, A2=>nx34775);
   max_calc_reg_comparator_third_inp1_7 : dff port map ( Q=>
      max_calc_comparator_third_inp1_7, QB=>nx30413, D=>nx21453, CLK=>clk);
   ix21454 : oai21 port map ( Y=>nx21453, A0=>nx30413, A1=>nx34775, B0=>
      nx30416);
   ix30417 : nand03 port map ( Y=>nx30416, A0=>label_5_output(7), A1=>
      nx35457, A2=>nx34775);
   ix30419 : aoi22 port map ( Y=>nx30418, A0=>nx30420, A1=>
      max_calc_comparator_third_inp1_6, B0=>nx12352, B1=>nx12530);
   max_calc_reg_comparator_third_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx30420, D=>nx21463, CLK=>clk);
   ix21464 : oai21 port map ( Y=>nx21463, A0=>nx30420, A1=>nx34775, B0=>
      nx30423);
   ix21474 : oai21 port map ( Y=>nx21473, A0=>nx30427, A1=>nx34775, B0=>
      nx30429);
   max_calc_reg_comparator_third_inp1_6 : dff port map ( Q=>
      max_calc_comparator_third_inp1_6, QB=>nx30427, D=>nx21473, CLK=>clk);
   ix12531 : oai22 port map ( Y=>nx12530, A0=>nx30433, A1=>nx30446, B0=>
      max_calc_comparator_third_inp2_5, B1=>nx30441);
   ix21484 : oai21 port map ( Y=>nx21483, A0=>nx30437, A1=>nx34777, B0=>
      nx30439);
   max_calc_reg_comparator_third_inp2_5 : dff port map ( Q=>
      max_calc_comparator_third_inp2_5, QB=>nx30437, D=>nx21483, CLK=>clk);
   ix30440 : nand03 port map ( Y=>nx30439, A0=>label_6_output(5), A1=>
      nx35457, A2=>nx34777);
   max_calc_reg_comparator_third_inp1_5 : dff port map ( Q=>
      max_calc_comparator_third_inp1_5, QB=>nx30441, D=>nx21493, CLK=>clk);
   ix21494 : oai21 port map ( Y=>nx21493, A0=>nx30441, A1=>nx34777, B0=>
      nx30444);
   ix30445 : nand03 port map ( Y=>nx30444, A0=>label_5_output(5), A1=>
      nx35459, A2=>nx34777);
   ix30447 : aoi22 port map ( Y=>nx30446, A0=>nx30448, A1=>
      max_calc_comparator_third_inp1_4, B0=>nx12396, B1=>nx12514);
   max_calc_reg_comparator_third_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx30448, D=>nx21503, CLK=>clk);
   ix21504 : oai21 port map ( Y=>nx21503, A0=>nx30448, A1=>nx34777, B0=>
      nx30451);
   ix21514 : oai21 port map ( Y=>nx21513, A0=>nx30455, A1=>nx34777, B0=>
      nx30457);
   max_calc_reg_comparator_third_inp1_4 : dff port map ( Q=>
      max_calc_comparator_third_inp1_4, QB=>nx30455, D=>nx21513, CLK=>clk);
   ix12515 : oai22 port map ( Y=>nx12514, A0=>nx30461, A1=>nx30474, B0=>
      max_calc_comparator_third_inp2_3, B1=>nx30469);
   ix21524 : oai21 port map ( Y=>nx21523, A0=>nx30465, A1=>nx34779, B0=>
      nx30467);
   max_calc_reg_comparator_third_inp2_3 : dff port map ( Q=>
      max_calc_comparator_third_inp2_3, QB=>nx30465, D=>nx21523, CLK=>clk);
   ix30468 : nand03 port map ( Y=>nx30467, A0=>label_6_output(3), A1=>
      nx35459, A2=>nx34779);
   max_calc_reg_comparator_third_inp1_3 : dff port map ( Q=>
      max_calc_comparator_third_inp1_3, QB=>nx30469, D=>nx21533, CLK=>clk);
   ix21534 : oai21 port map ( Y=>nx21533, A0=>nx30469, A1=>nx34779, B0=>
      nx30472);
   ix30473 : nand03 port map ( Y=>nx30472, A0=>label_5_output(3), A1=>
      nx35459, A2=>nx34779);
   ix30475 : aoi22 port map ( Y=>nx30474, A0=>nx30476, A1=>
      max_calc_comparator_third_inp1_2, B0=>nx12440, B1=>nx12498);
   max_calc_reg_comparator_third_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx30476, D=>nx21543, CLK=>clk);
   ix21544 : oai21 port map ( Y=>nx21543, A0=>nx30476, A1=>nx34779, B0=>
      nx30479);
   ix21554 : oai21 port map ( Y=>nx21553, A0=>nx30483, A1=>nx34781, B0=>
      nx30485);
   max_calc_reg_comparator_third_inp1_2 : dff port map ( Q=>
      max_calc_comparator_third_inp1_2, QB=>nx30483, D=>nx21553, CLK=>clk);
   ix12499 : oai21 port map ( Y=>nx12498, A0=>
      max_calc_comparator_third_inp2_1, A1=>nx30495, B0=>nx30500);
   ix21564 : oai21 port map ( Y=>nx21563, A0=>nx30491, A1=>nx34781, B0=>
      nx30493);
   max_calc_reg_comparator_third_inp2_1 : dff port map ( Q=>
      max_calc_comparator_third_inp2_1, QB=>nx30491, D=>nx21563, CLK=>clk);
   ix30494 : nand03 port map ( Y=>nx30493, A0=>label_6_output(1), A1=>
      nx35461, A2=>nx34781);
   max_calc_reg_comparator_third_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx30495, D=>nx21573, CLK=>clk);
   ix21574 : oai21 port map ( Y=>nx21573, A0=>nx30495, A1=>nx34781, B0=>
      nx30498);
   ix30499 : nand03 port map ( Y=>nx30498, A0=>label_5_output(1), A1=>
      nx35461, A2=>nx34781);
   ix30501 : oai21 port map ( Y=>nx30500, A0=>nx29502, A1=>
      max_calc_comparator_third_inp1_0, B0=>nx12462);
   ix21624 : oai21 port map ( Y=>nx21623, A0=>nx30506, A1=>nx34781, B0=>
      nx30508);
   max_calc_reg_comparator_third_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx30506, D=>nx21623, CLK=>clk);
   ix30509 : nand03 port map ( Y=>nx30508, A0=>label_6_output(15), A1=>
      nx35461, A2=>nx34783);
   labelsregfile_label6_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_6_output(15), QB=>OPEN, D=>nx21613, CLK=>clk, R=>rst);
   lat_label_6_input_15 : latch port map ( Q=>label_6_input_15, D=>nx12624, 
      CLK=>nx34529);
   reg_label_6_input_state_machine_15 : dffr port map ( Q=>
      label_6_input_state_machine_15, QB=>OPEN, D=>nx21603, CLK=>clk, R=>rst
   );
   ix12621 : xnor2 port map ( Y=>nx12620, A0=>nx12616, A1=>nx30519);
   ix12617 : oai22 port map ( Y=>nx12616, A0=>nx29955, A1=>nx30127, B0=>
      nx30129, B1=>nx29923);
   ix21654 : oai21 port map ( Y=>nx21653, A0=>nx30524, A1=>nx34783, B0=>
      nx30526);
   max_calc_reg_comparator_third_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx30524, D=>nx21653, CLK=>clk);
   ix30527 : nand03 port map ( Y=>nx30526, A0=>label_5_output(15), A1=>
      nx35461, A2=>nx34783);
   labelsregfile_label5_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_5_output(15), QB=>OPEN, D=>nx21643, CLK=>clk, R=>rst);
   lat_label_5_input_15 : latch port map ( Q=>label_5_input_15, D=>nx12666, 
      CLK=>nx34529);
   reg_label_5_input_state_machine_15 : dffr port map ( Q=>
      label_5_input_state_machine_15, QB=>OPEN, D=>nx21633, CLK=>clk, R=>rst
   );
   ix12663 : xnor2 port map ( Y=>nx12662, A0=>nx12658, A1=>nx30537);
   ix12659 : oai22 port map ( Y=>nx12658, A0=>nx30144, A1=>nx30316, B0=>
      nx30318, B1=>nx29482);
   max_calc_reg_ans3_0 : dff port map ( Q=>max_calc_ans3_0, QB=>OPEN, D=>
      nx24263, CLK=>clk);
   ix24254 : oai21 port map ( Y=>nx24253, A0=>nx30546, A1=>nx34783, B0=>
      nx30548);
   max_calc_reg_comparator_second_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx30546, D=>nx24253, CLK=>clk);
   ix30549 : nand03 port map ( Y=>nx30548, A0=>nx35175, A1=>nx16896, A2=>
      nx34801);
   labelsregfile_label4_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_4_output(0), QB=>OPEN, D=>nx14673, CLK=>clk, R=>rst);
   lat_label_4_input_0 : latch port map ( Q=>label_4_input_0, D=>nx1744, CLK
      =>nx34529);
   ix1745 : oai21 port map ( Y=>nx1744, A0=>nx30555, A1=>nx34429, B0=>
      nx30559);
   reg_label_4_input_state_machine_0 : dffr port map ( Q=>
      label_4_input_state_machine_0, QB=>nx30555, D=>nx14663, CLK=>clk, R=>
      rst);
   ix30560 : oai21 port map ( Y=>nx30559, A0=>nx35719, A1=>label_4_output(0), 
      B0=>nx1732);
   booth_booth_integrtaion_3_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_1, QB=>OPEN, D=>nx14643, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_2, QB=>nx30980, D=>nx14633, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_3, QB=>OPEN, D=>nx14623, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_4, QB=>nx30978, D=>nx14613, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_5, QB=>OPEN, D=>nx14603, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_6, QB=>nx30976, D=>nx14593, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_7, QB=>OPEN, D=>nx14583, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_8, QB=>nx30974, D=>nx14573, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_9, QB=>OPEN, D=>nx14563, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_10, QB=>nx30972, D=>nx14553, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_11, QB=>OPEN, D=>nx14543, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_12, QB=>nx30970, D=>nx14533, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_13, QB=>OPEN, D=>nx14523, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_14, QB=>nx30968, D=>nx14513, CLK=>clk, 
      R=>rst);
   ix30609 : aoi22 port map ( Y=>nx30608, A0=>mdr_data_out(15), A1=>nx34571, 
      B0=>nx1530, B1=>nx1536);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_reg_output_0, QB=>OPEN, 
      D=>nx14153, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_0, QB=>OPEN, D=>nx14139, CLK
      =>clk, S=>nx34487);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_reg_output_9, QB=>OPEN, 
      D=>nx14333, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_9, QB=>OPEN, D=>nx14323, CLK
      =>clk, R=>nx34487);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_8, QB=>OPEN, 
      D=>nx14313, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_8, QB=>OPEN, D=>nx14303, CLK
      =>clk, R=>nx34487);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_7, QB=>OPEN, 
      D=>nx14293, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_7, QB=>OPEN, D=>nx14283, CLK
      =>clk, R=>nx34485);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_6, QB=>OPEN, 
      D=>nx14273, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_6, QB=>OPEN, D=>nx14263, CLK
      =>clk, R=>nx34485);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_5, QB=>OPEN, 
      D=>nx14253, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_5, QB=>OPEN, D=>nx14243, CLK
      =>clk, R=>nx34485);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_4, QB=>OPEN, 
      D=>nx14233, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_4, QB=>OPEN, D=>nx14223, CLK
      =>clk, R=>nx34485);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_3, QB=>OPEN, 
      D=>nx14213, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_3, QB=>OPEN, D=>nx14203, CLK
      =>clk, R=>nx34485);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_2, QB=>OPEN, 
      D=>nx14193, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_2, QB=>OPEN, D=>nx14183, CLK
      =>clk, R=>nx34485);
   booth_booth_integrtaion_3_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_3_shift_Reg_output_1, QB=>OPEN, 
      D=>nx14173, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_3_shift_Reg_count_1, QB=>OPEN, D=>nx14163, CLK
      =>clk, R=>nx34483);
   ix14134 : nand02 port map ( Y=>nx14133, A0=>nx35831, A1=>nx34557);
   booth_booth_integrtaion_3_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx30655, D=>nx14133, CLK=>clk, S=>nx34485);
   ix1531 : nand02 port map ( Y=>nx1530, A0=>nx30676, A1=>nx30688);
   ix30677 : oai21 port map ( Y=>nx30676, A0=>nx34585, A1=>nx34579, B0=>
      mdr_data_out(64));
   ix14344 : oai21 port map ( Y=>nx14343, A0=>nx30681, A1=>nx35499, B0=>
      nx30683);
   booth_booth_integrtaion_3_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx30681, D=>nx14343, CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx30685, D=>nx14653, CLK=>clk, R=>rst);
   ix30693 : xnor2 port map ( Y=>nx30692, A0=>nx1000, A1=>nx12913);
   ix14484 : oai21 port map ( Y=>nx14483, A0=>nx30698, A1=>nx35499, B0=>
      nx30700);
   booth_booth_integrtaion_3_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_17, QB=>nx30698, D=>nx14483, 
      CLK=>clk, R=>rst);
   ix30701 : nand03 port map ( Y=>nx30700, A0=>nx35507, A1=>nx1508, A2=>
      nx36147);
   ix1509 : xnor2 port map ( Y=>nx1508, A0=>nx30703, A1=>nx12915);
   ix30704 : aoi22 port map ( Y=>nx30703, A0=>
      booth_booth_integrtaion_3_booth_output_17, A1=>nx1024, B0=>nx1000, B1
      =>nx12913);
   ix1009 : nand02 port map ( Y=>nx1008, A0=>mdr_data_out(65), A1=>
      mdr_data_out(64));
   ix30708 : or02 port map ( Y=>nx30707, A0=>mdr_data_out(64), A1=>
      mdr_data_out(65));
   ix30714 : xnor2 port map ( Y=>nx30713, A0=>nx1052, A1=>nx12917);
   ix1053 : oai22 port map ( Y=>nx1052, A0=>nx30703, A1=>nx30716, B0=>
      nx30723, B1=>nx35511);
   ix30719 : aoi32 port map ( Y=>nx30718, A0=>nx1034, A1=>nx34585, A2=>
      nx30721, B0=>mdr_data_out(66), B1=>nx34579);
   ix1035 : oai21 port map ( Y=>nx1034, A0=>mdr_data_out(64), A1=>
      mdr_data_out(65), B0=>mdr_data_out(66));
   booth_booth_integrtaion_3_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_18, QB=>nx30723, D=>nx14473, 
      CLK=>clk, R=>rst);
   ix14464 : oai21 port map ( Y=>nx14463, A0=>nx30728, A1=>nx35499, B0=>
      nx30730);
   booth_booth_integrtaion_3_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_19, QB=>nx30728, D=>nx14463, 
      CLK=>clk, R=>rst);
   ix30731 : nand03 port map ( Y=>nx30730, A0=>nx35507, A1=>nx1484, A2=>
      nx36147);
   ix1485 : xnor2 port map ( Y=>nx1484, A0=>nx30733, A1=>nx12919);
   ix30734 : aoi22 port map ( Y=>nx30733, A0=>
      booth_booth_integrtaion_3_booth_output_19, A1=>nx1072, B0=>nx1052, B1
      =>nx12917);
   ix30737 : nor02ii port map ( Y=>nx30736, A0=>nx1038, A1=>mdr_data_out(67)
   );
   ix1039 : nor03_2x port map ( Y=>nx1038, A0=>mdr_data_out(66), A1=>
      mdr_data_out(64), A2=>mdr_data_out(65));
   ix1063 : nor04 port map ( Y=>nx1062, A0=>mdr_data_out(67), A1=>
      mdr_data_out(66), A2=>mdr_data_out(64), A3=>mdr_data_out(65));
   ix30751 : xnor2 port map ( Y=>nx30750, A0=>nx1100, A1=>nx12921);
   ix1101 : oai22 port map ( Y=>nx1100, A0=>nx30733, A1=>nx30753, B0=>
      nx30762, B1=>nx35513);
   ix30756 : aoi32 port map ( Y=>nx30755, A0=>nx1082, A1=>nx34585, A2=>
      nx30760, B0=>mdr_data_out(68), B1=>nx34579);
   ix1083 : nand02 port map ( Y=>nx1082, A0=>nx30758, A1=>mdr_data_out(68));
   booth_booth_integrtaion_3_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_20, QB=>nx30762, D=>nx14453, 
      CLK=>clk, R=>rst);
   ix14444 : oai21 port map ( Y=>nx14443, A0=>nx30767, A1=>nx35499, B0=>
      nx30769);
   booth_booth_integrtaion_3_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_21, QB=>nx30767, D=>nx14443, 
      CLK=>clk, R=>rst);
   ix30770 : nand03 port map ( Y=>nx30769, A0=>nx35507, A1=>nx1460, A2=>
      nx36147);
   ix1461 : xnor2 port map ( Y=>nx1460, A0=>nx30772, A1=>nx12922);
   ix30773 : aoi22 port map ( Y=>nx30772, A0=>
      booth_booth_integrtaion_3_booth_output_21, A1=>nx1120, B0=>nx1100, B1
      =>nx12921);
   ix30776 : nor02ii port map ( Y=>nx30775, A0=>nx1086, A1=>mdr_data_out(69)
   );
   ix1087 : nor02ii port map ( Y=>nx1086, A0=>mdr_data_out(68), A1=>nx1062);
   ix1111 : nor02ii port map ( Y=>nx1110, A0=>mdr_data_out(69), A1=>nx1086);
   ix30786 : xnor2 port map ( Y=>nx30785, A0=>nx1148, A1=>nx12923);
   ix1149 : oai22 port map ( Y=>nx1148, A0=>nx30772, A1=>nx30788, B0=>
      nx30797, B1=>nx35515);
   ix30791 : aoi32 port map ( Y=>nx30790, A0=>nx1130, A1=>nx34585, A2=>
      nx30795, B0=>mdr_data_out(70), B1=>nx34579);
   ix1131 : nand02 port map ( Y=>nx1130, A0=>nx30793, A1=>mdr_data_out(70));
   booth_booth_integrtaion_3_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_22, QB=>nx30797, D=>nx14433, 
      CLK=>clk, R=>rst);
   ix14424 : oai21 port map ( Y=>nx14423, A0=>nx30802, A1=>nx35499, B0=>
      nx30804);
   booth_booth_integrtaion_3_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_23, QB=>nx30802, D=>nx14423, 
      CLK=>clk, R=>rst);
   ix30805 : nand03 port map ( Y=>nx30804, A0=>nx35507, A1=>nx1436, A2=>
      nx35501);
   ix1437 : xnor2 port map ( Y=>nx1436, A0=>nx30807, A1=>nx12925);
   ix30808 : aoi22 port map ( Y=>nx30807, A0=>
      booth_booth_integrtaion_3_booth_output_23, A1=>nx1168, B0=>nx1148, B1
      =>nx12923);
   ix30811 : nor02ii port map ( Y=>nx30810, A0=>nx1134, A1=>mdr_data_out(71)
   );
   ix1135 : nor02ii port map ( Y=>nx1134, A0=>mdr_data_out(70), A1=>nx1110);
   ix1159 : nor02ii port map ( Y=>nx1158, A0=>mdr_data_out(71), A1=>nx1134);
   ix30821 : xnor2 port map ( Y=>nx30820, A0=>nx1196, A1=>nx12927);
   ix1197 : oai22 port map ( Y=>nx1196, A0=>nx30807, A1=>nx30823, B0=>
      nx30832, B1=>nx35517);
   ix30826 : aoi32 port map ( Y=>nx30825, A0=>nx1178, A1=>nx34585, A2=>
      nx30830, B0=>mdr_data_out(72), B1=>nx34579);
   ix1179 : nand02 port map ( Y=>nx1178, A0=>nx30828, A1=>mdr_data_out(72));
   booth_booth_integrtaion_3_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_24, QB=>nx30832, D=>nx14413, 
      CLK=>clk, R=>rst);
   ix14404 : oai21 port map ( Y=>nx14403, A0=>nx30837, A1=>nx35501, B0=>
      nx30839);
   booth_booth_integrtaion_3_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_25, QB=>nx30837, D=>nx14403, 
      CLK=>clk, R=>rst);
   ix30840 : nand03 port map ( Y=>nx30839, A0=>nx35507, A1=>nx1412, A2=>
      nx35501);
   ix1413 : xnor2 port map ( Y=>nx1412, A0=>nx30842, A1=>nx12929);
   ix30843 : aoi22 port map ( Y=>nx30842, A0=>
      booth_booth_integrtaion_3_booth_output_25, A1=>nx1216, B0=>nx1196, B1
      =>nx12927);
   ix30846 : nor02ii port map ( Y=>nx30845, A0=>nx1182, A1=>mdr_data_out(73)
   );
   ix1183 : nor02ii port map ( Y=>nx1182, A0=>mdr_data_out(72), A1=>nx1158);
   ix1207 : nor02ii port map ( Y=>nx1206, A0=>mdr_data_out(73), A1=>nx1182);
   ix30856 : xnor2 port map ( Y=>nx30855, A0=>nx1244, A1=>nx12930);
   ix1245 : oai22 port map ( Y=>nx1244, A0=>nx30842, A1=>nx30858, B0=>
      nx30867, B1=>nx35519);
   ix30861 : aoi32 port map ( Y=>nx30860, A0=>nx1226, A1=>nx34585, A2=>
      nx30865, B0=>mdr_data_out(74), B1=>nx34579);
   ix1227 : nand02 port map ( Y=>nx1226, A0=>nx30863, A1=>mdr_data_out(74));
   booth_booth_integrtaion_3_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_26, QB=>nx30867, D=>nx14393, 
      CLK=>clk, R=>rst);
   ix14384 : oai21 port map ( Y=>nx14383, A0=>nx30872, A1=>nx35501, B0=>
      nx30874);
   booth_booth_integrtaion_3_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_27, QB=>nx30872, D=>nx14383, 
      CLK=>clk, R=>rst);
   ix30875 : nand03 port map ( Y=>nx30874, A0=>nx35507, A1=>nx1388, A2=>
      nx35501);
   ix1389 : xnor2 port map ( Y=>nx1388, A0=>nx30877, A1=>nx12931);
   ix30878 : aoi22 port map ( Y=>nx30877, A0=>
      booth_booth_integrtaion_3_booth_output_27, A1=>nx1264, B0=>nx1244, B1
      =>nx12930);
   ix30881 : nor02ii port map ( Y=>nx30880, A0=>nx1230, A1=>mdr_data_out(75)
   );
   ix1231 : nor02ii port map ( Y=>nx1230, A0=>mdr_data_out(74), A1=>nx1206);
   ix1255 : nor02ii port map ( Y=>nx1254, A0=>mdr_data_out(75), A1=>nx1230);
   ix30891 : xnor2 port map ( Y=>nx30890, A0=>nx1292, A1=>nx12933);
   ix1293 : oai22 port map ( Y=>nx1292, A0=>nx30877, A1=>nx30893, B0=>
      nx30902, B1=>nx35521);
   ix30896 : aoi32 port map ( Y=>nx30895, A0=>nx1274, A1=>nx34585, A2=>
      nx30900, B0=>mdr_data_out(76), B1=>nx34579);
   ix1275 : nand02 port map ( Y=>nx1274, A0=>nx30898, A1=>mdr_data_out(76));
   booth_booth_integrtaion_3_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_28, QB=>nx30902, D=>nx14373, 
      CLK=>clk, R=>rst);
   ix14364 : oai21 port map ( Y=>nx14363, A0=>nx30907, A1=>nx35501, B0=>
      nx30909);
   booth_booth_integrtaion_3_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_29, QB=>nx30907, D=>nx14363, 
      CLK=>clk, R=>rst);
   ix30910 : nand03 port map ( Y=>nx30909, A0=>nx36155, A1=>nx1364, A2=>
      nx35501);
   ix1365 : xnor2 port map ( Y=>nx1364, A0=>nx30912, A1=>nx12935);
   ix30913 : aoi22 port map ( Y=>nx30912, A0=>
      booth_booth_integrtaion_3_booth_output_29, A1=>nx1312, B0=>nx1292, B1
      =>nx12933);
   ix30916 : nor02ii port map ( Y=>nx30915, A0=>nx1278, A1=>mdr_data_out(77)
   );
   ix1279 : nor02ii port map ( Y=>nx1278, A0=>mdr_data_out(76), A1=>nx1254);
   ix1303 : nor02ii port map ( Y=>nx1302, A0=>mdr_data_out(77), A1=>nx1278);
   ix30926 : xnor2 port map ( Y=>nx30925, A0=>nx1340, A1=>nx1350);
   ix1341 : oai22 port map ( Y=>nx1340, A0=>nx30912, A1=>nx30928, B0=>
      nx30937, B1=>nx35523);
   ix30931 : aoi32 port map ( Y=>nx30930, A0=>nx1322, A1=>nx34587, A2=>
      nx30935, B0=>mdr_data_out(78), B1=>nx34581);
   ix1323 : nand02 port map ( Y=>nx1322, A0=>nx30933, A1=>mdr_data_out(78));
   booth_booth_integrtaion_3_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_31, QB=>nx30937, D=>nx14353, 
      CLK=>clk, R=>rst);
   ix30941 : aoi22 port map ( Y=>nx30940, A0=>mdr_data_out(79), A1=>nx34581, 
      B0=>nx34587, B1=>nx1342);
   ix1343 : xnor2 port map ( Y=>nx1342, A0=>mdr_data_out(79), A1=>nx1326);
   ix1327 : nor02ii port map ( Y=>nx1326, A0=>mdr_data_out(78), A1=>nx1302);
   ix30945 : aoi32 port map ( Y=>nx30944, A0=>nx1298, A1=>nx34587, A2=>
      nx30933, B0=>mdr_data_out(77), B1=>nx34581);
   ix30948 : aoi32 port map ( Y=>nx30947, A0=>nx1250, A1=>nx34587, A2=>
      nx30898, B0=>mdr_data_out(75), B1=>nx34581);
   ix30951 : aoi32 port map ( Y=>nx30950, A0=>nx1202, A1=>nx34587, A2=>
      nx30863, B0=>mdr_data_out(73), B1=>nx34581);
   ix30954 : aoi32 port map ( Y=>nx30953, A0=>nx1154, A1=>nx34587, A2=>
      nx30828, B0=>mdr_data_out(71), B1=>nx34581);
   ix30957 : aoi32 port map ( Y=>nx30956, A0=>nx1106, A1=>nx34587, A2=>
      nx30793, B0=>mdr_data_out(69), B1=>nx34581);
   ix30960 : aoi32 port map ( Y=>nx30959, A0=>nx1058, A1=>nx994, A2=>nx30758, 
      B0=>mdr_data_out(67), B1=>nx34583);
   ix30963 : aoi32 port map ( Y=>nx30962, A0=>nx1008, A1=>nx994, A2=>nx30707, 
      B0=>mdr_data_out(65), B1=>nx34583);
   booth_booth_integrtaion_3_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_3_booth_output_16, QB=>nx30688, D=>nx14493, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_3_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_3_15, QB=>nx30966, D=>nx14503, CLK=>clk, 
      R=>rst);
   ix1733 : aoi21 port map ( Y=>nx1732, A0=>label_4_output(0), A1=>nx35719, 
      B0=>nx35919);
   ix23634 : oai21 port map ( Y=>nx23633, A0=>nx30990, A1=>nx34783, B0=>
      nx30992);
   max_calc_reg_comparator_fourth_inp1_0 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_0, QB=>nx30990, D=>nx23633, CLK=>clk);
   ix30993 : nand03 port map ( Y=>nx30992, A0=>label_7_output(0), A1=>
      nx35461, A2=>nx34783);
   labelsregfile_label7_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_7_output(0), QB=>OPEN, D=>nx22233, CLK=>clk, R=>rst);
   lat_label_7_input_0 : latch port map ( Q=>label_7_input_0, D=>nx13586, 
      CLK=>nx34529);
   ix13587 : oai21 port map ( Y=>nx13586, A0=>nx30998, A1=>nx34429, B0=>
      nx31002);
   reg_label_7_input_state_machine_0 : dffr port map ( Q=>
      label_7_input_state_machine_0, QB=>nx30998, D=>nx22223, CLK=>clk, R=>
      rst);
   ix31003 : oai21 port map ( Y=>nx31002, A0=>nx35771, A1=>label_7_output(0), 
      B0=>nx13574);
   booth_booth_integrtaion_6_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_1, QB=>OPEN, D=>nx22203, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_2, QB=>nx31423, D=>nx22193, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_3, QB=>OPEN, D=>nx22183, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_4, QB=>nx31421, D=>nx22173, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_5, QB=>OPEN, D=>nx22163, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_6, QB=>nx31419, D=>nx22153, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_7, QB=>OPEN, D=>nx22143, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_8, QB=>nx31417, D=>nx22133, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_9, QB=>OPEN, D=>nx22123, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_10, QB=>nx31415, D=>nx22113, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_11, QB=>OPEN, D=>nx22103, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_12, QB=>nx31413, D=>nx22093, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_13, QB=>OPEN, D=>nx22083, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_14, QB=>nx31411, D=>nx22073, CLK=>clk, 
      R=>rst);
   ix31052 : aoi22 port map ( Y=>nx31051, A0=>mdr_data_out(15), A1=>nx35011, 
      B0=>nx13372, B1=>nx13378);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_reg_output_0, QB=>OPEN, 
      D=>nx21713, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_0, QB=>OPEN, D=>nx21699, CLK
      =>clk, S=>nx34489);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_reg_output_9, QB=>OPEN, 
      D=>nx21893, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_9, QB=>OPEN, D=>nx21883, CLK
      =>clk, R=>nx34489);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_8, QB=>OPEN, 
      D=>nx21873, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_8, QB=>OPEN, D=>nx21863, CLK
      =>clk, R=>nx34489);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_7, QB=>OPEN, 
      D=>nx21853, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_7, QB=>OPEN, D=>nx21843, CLK
      =>clk, R=>nx34489);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_6, QB=>OPEN, 
      D=>nx21833, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_6, QB=>OPEN, D=>nx21823, CLK
      =>clk, R=>nx34489);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_5, QB=>OPEN, 
      D=>nx21813, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_5, QB=>OPEN, D=>nx21803, CLK
      =>clk, R=>nx34489);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_4, QB=>OPEN, 
      D=>nx21793, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_4, QB=>OPEN, D=>nx21783, CLK
      =>clk, R=>nx34489);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_3, QB=>OPEN, 
      D=>nx21773, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_3, QB=>OPEN, D=>nx21763, CLK
      =>clk, R=>nx34487);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_2, QB=>OPEN, 
      D=>nx21753, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_2, QB=>OPEN, D=>nx21743, CLK
      =>clk, R=>nx34487);
   booth_booth_integrtaion_6_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_6_shift_Reg_output_1, QB=>OPEN, 
      D=>nx21733, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_6_shift_Reg_count_1, QB=>OPEN, D=>nx21723, CLK
      =>clk, R=>nx34487);
   ix21694 : nand02 port map ( Y=>nx21693, A0=>nx35835, A1=>nx34997);
   booth_booth_integrtaion_6_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx31098, D=>nx21693, CLK=>clk, S=>nx34487);
   ix13373 : nand02 port map ( Y=>nx13372, A0=>nx31119, A1=>nx31131);
   ix31120 : oai21 port map ( Y=>nx31119, A0=>nx35025, A1=>nx35019, B0=>
      mdr_data_out(112));
   ix21904 : oai21 port map ( Y=>nx21903, A0=>nx31124, A1=>nx35525, B0=>
      nx31126);
   booth_booth_integrtaion_6_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx31124, D=>nx21903, CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx31128, D=>nx22213, CLK=>clk, R=>rst);
   ix31136 : xnor2 port map ( Y=>nx31135, A0=>nx12842, A1=>nx13296);
   ix22044 : oai21 port map ( Y=>nx22043, A0=>nx31141, A1=>nx35525, B0=>
      nx31143);
   booth_booth_integrtaion_6_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_17, QB=>nx31141, D=>nx22043, 
      CLK=>clk, R=>rst);
   ix31144 : nand03 port map ( Y=>nx31143, A0=>nx35533, A1=>nx13350, A2=>
      nx36163);
   ix13351 : xnor2 port map ( Y=>nx13350, A0=>nx31146, A1=>nx13297);
   ix31147 : aoi22 port map ( Y=>nx31146, A0=>
      booth_booth_integrtaion_6_booth_output_17, A1=>nx12866, B0=>nx12842, 
      B1=>nx13296);
   ix12851 : nand02 port map ( Y=>nx12850, A0=>mdr_data_out(113), A1=>
      mdr_data_out(112));
   ix31151 : or02 port map ( Y=>nx31150, A0=>mdr_data_out(112), A1=>
      mdr_data_out(113));
   ix31157 : xnor2 port map ( Y=>nx31156, A0=>nx12894, A1=>nx13298);
   ix12895 : oai22 port map ( Y=>nx12894, A0=>nx31146, A1=>nx31159, B0=>
      nx31166, B1=>nx35537);
   ix31162 : aoi32 port map ( Y=>nx31161, A0=>nx12876, A1=>nx35025, A2=>
      nx31164, B0=>mdr_data_out(114), B1=>nx35019);
   ix12877 : oai21 port map ( Y=>nx12876, A0=>mdr_data_out(112), A1=>
      mdr_data_out(113), B0=>mdr_data_out(114));
   booth_booth_integrtaion_6_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_18, QB=>nx31166, D=>nx22033, 
      CLK=>clk, R=>rst);
   ix22024 : oai21 port map ( Y=>nx22023, A0=>nx31171, A1=>nx35525, B0=>
      nx31173);
   booth_booth_integrtaion_6_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_19, QB=>nx31171, D=>nx22023, 
      CLK=>clk, R=>rst);
   ix31174 : nand03 port map ( Y=>nx31173, A0=>nx35533, A1=>nx13326, A2=>
      nx36163);
   ix13327 : xnor2 port map ( Y=>nx13326, A0=>nx31176, A1=>nx13299);
   ix31177 : aoi22 port map ( Y=>nx31176, A0=>
      booth_booth_integrtaion_6_booth_output_19, A1=>nx12914, B0=>nx12894, 
      B1=>nx13298);
   ix31180 : nor02ii port map ( Y=>nx31179, A0=>nx12880, A1=>
      mdr_data_out(115));
   ix12881 : nor03_2x port map ( Y=>nx12880, A0=>mdr_data_out(114), A1=>
      mdr_data_out(112), A2=>mdr_data_out(113));
   ix12905 : nor04 port map ( Y=>nx12904, A0=>mdr_data_out(115), A1=>
      mdr_data_out(114), A2=>mdr_data_out(112), A3=>mdr_data_out(113));
   ix31194 : xnor2 port map ( Y=>nx31193, A0=>nx12942, A1=>nx13300);
   ix12943 : oai22 port map ( Y=>nx12942, A0=>nx31176, A1=>nx31196, B0=>
      nx31205, B1=>nx35539);
   ix31199 : aoi32 port map ( Y=>nx31198, A0=>nx12924, A1=>nx35025, A2=>
      nx31203, B0=>mdr_data_out(116), B1=>nx35019);
   ix12925 : nand02 port map ( Y=>nx12924, A0=>nx31201, A1=>
      mdr_data_out(116));
   booth_booth_integrtaion_6_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_20, QB=>nx31205, D=>nx22013, 
      CLK=>clk, R=>rst);
   ix22004 : oai21 port map ( Y=>nx22003, A0=>nx31210, A1=>nx35525, B0=>
      nx31212);
   booth_booth_integrtaion_6_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_21, QB=>nx31210, D=>nx22003, 
      CLK=>clk, R=>rst);
   ix31213 : nand03 port map ( Y=>nx31212, A0=>nx35533, A1=>nx13302, A2=>
      nx36163);
   ix13303 : xnor2 port map ( Y=>nx13302, A0=>nx31215, A1=>nx13301);
   ix31216 : aoi22 port map ( Y=>nx31215, A0=>
      booth_booth_integrtaion_6_booth_output_21, A1=>nx12962, B0=>nx12942, 
      B1=>nx13300);
   ix31219 : nor02ii port map ( Y=>nx31218, A0=>nx12928, A1=>
      mdr_data_out(117));
   ix12929 : nor02ii port map ( Y=>nx12928, A0=>mdr_data_out(116), A1=>
      nx12904);
   ix12953 : nor02ii port map ( Y=>nx12952, A0=>mdr_data_out(117), A1=>
      nx12928);
   ix31229 : xnor2 port map ( Y=>nx31228, A0=>nx12990, A1=>nx13303);
   ix12991 : oai22 port map ( Y=>nx12990, A0=>nx31215, A1=>nx31231, B0=>
      nx31240, B1=>nx35541);
   ix31234 : aoi32 port map ( Y=>nx31233, A0=>nx12972, A1=>nx35025, A2=>
      nx31238, B0=>mdr_data_out(118), B1=>nx35019);
   ix12973 : nand02 port map ( Y=>nx12972, A0=>nx31236, A1=>
      mdr_data_out(118));
   booth_booth_integrtaion_6_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_22, QB=>nx31240, D=>nx21993, 
      CLK=>clk, R=>rst);
   ix21984 : oai21 port map ( Y=>nx21983, A0=>nx31245, A1=>nx35525, B0=>
      nx31247);
   booth_booth_integrtaion_6_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_23, QB=>nx31245, D=>nx21983, 
      CLK=>clk, R=>rst);
   ix31248 : nand03 port map ( Y=>nx31247, A0=>nx35533, A1=>nx13278, A2=>
      nx35527);
   ix13279 : xnor2 port map ( Y=>nx13278, A0=>nx31250, A1=>nx13305);
   ix31251 : aoi22 port map ( Y=>nx31250, A0=>
      booth_booth_integrtaion_6_booth_output_23, A1=>nx13010, B0=>nx12990, 
      B1=>nx13303);
   ix31254 : nor02ii port map ( Y=>nx31253, A0=>nx12976, A1=>
      mdr_data_out(119));
   ix12977 : nor02ii port map ( Y=>nx12976, A0=>mdr_data_out(118), A1=>
      nx12952);
   ix13001 : nor02ii port map ( Y=>nx13000, A0=>mdr_data_out(119), A1=>
      nx12976);
   ix31264 : xnor2 port map ( Y=>nx31263, A0=>nx13038, A1=>nx13307);
   ix13039 : oai22 port map ( Y=>nx13038, A0=>nx31250, A1=>nx31266, B0=>
      nx31275, B1=>nx35543);
   ix31269 : aoi32 port map ( Y=>nx31268, A0=>nx13020, A1=>nx35025, A2=>
      nx31273, B0=>mdr_data_out(120), B1=>nx35019);
   ix13021 : nand02 port map ( Y=>nx13020, A0=>nx31271, A1=>
      mdr_data_out(120));
   booth_booth_integrtaion_6_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_24, QB=>nx31275, D=>nx21973, 
      CLK=>clk, R=>rst);
   ix21964 : oai21 port map ( Y=>nx21963, A0=>nx31280, A1=>nx35527, B0=>
      nx31282);
   booth_booth_integrtaion_6_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_25, QB=>nx31280, D=>nx21963, 
      CLK=>clk, R=>rst);
   ix31283 : nand03 port map ( Y=>nx31282, A0=>nx35533, A1=>nx13254, A2=>
      nx35527);
   ix13255 : xnor2 port map ( Y=>nx13254, A0=>nx31285, A1=>nx13308);
   ix31286 : aoi22 port map ( Y=>nx31285, A0=>
      booth_booth_integrtaion_6_booth_output_25, A1=>nx13058, B0=>nx13038, 
      B1=>nx13307);
   ix31289 : nor02ii port map ( Y=>nx31288, A0=>nx13024, A1=>
      mdr_data_out(121));
   ix13025 : nor02ii port map ( Y=>nx13024, A0=>mdr_data_out(120), A1=>
      nx13000);
   ix13049 : nor02ii port map ( Y=>nx13048, A0=>mdr_data_out(121), A1=>
      nx13024);
   ix31299 : xnor2 port map ( Y=>nx31298, A0=>nx13086, A1=>nx13309);
   ix13087 : oai22 port map ( Y=>nx13086, A0=>nx31285, A1=>nx31301, B0=>
      nx31310, B1=>nx35545);
   ix31304 : aoi32 port map ( Y=>nx31303, A0=>nx13068, A1=>nx35025, A2=>
      nx31308, B0=>mdr_data_out(122), B1=>nx35019);
   ix13069 : nand02 port map ( Y=>nx13068, A0=>nx31306, A1=>
      mdr_data_out(122));
   booth_booth_integrtaion_6_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_26, QB=>nx31310, D=>nx21953, 
      CLK=>clk, R=>rst);
   ix21944 : oai21 port map ( Y=>nx21943, A0=>nx31315, A1=>nx35527, B0=>
      nx31317);
   booth_booth_integrtaion_6_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_27, QB=>nx31315, D=>nx21943, 
      CLK=>clk, R=>rst);
   ix31318 : nand03 port map ( Y=>nx31317, A0=>nx35533, A1=>nx13230, A2=>
      nx35527);
   ix13231 : xnor2 port map ( Y=>nx13230, A0=>nx31320, A1=>nx13310);
   ix31321 : aoi22 port map ( Y=>nx31320, A0=>
      booth_booth_integrtaion_6_booth_output_27, A1=>nx13106, B0=>nx13086, 
      B1=>nx13309);
   ix31324 : nor02ii port map ( Y=>nx31323, A0=>nx13072, A1=>
      mdr_data_out(123));
   ix13073 : nor02ii port map ( Y=>nx13072, A0=>mdr_data_out(122), A1=>
      nx13048);
   ix13097 : nor02ii port map ( Y=>nx13096, A0=>mdr_data_out(123), A1=>
      nx13072);
   ix31334 : xnor2 port map ( Y=>nx31333, A0=>nx13134, A1=>nx13311);
   ix13135 : oai22 port map ( Y=>nx13134, A0=>nx31320, A1=>nx31336, B0=>
      nx31345, B1=>nx35547);
   ix31339 : aoi32 port map ( Y=>nx31338, A0=>nx13116, A1=>nx35025, A2=>
      nx31343, B0=>mdr_data_out(124), B1=>nx35019);
   ix13117 : nand02 port map ( Y=>nx13116, A0=>nx31341, A1=>
      mdr_data_out(124));
   booth_booth_integrtaion_6_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_28, QB=>nx31345, D=>nx21933, 
      CLK=>clk, R=>rst);
   ix21924 : oai21 port map ( Y=>nx21923, A0=>nx31350, A1=>nx35527, B0=>
      nx31352);
   booth_booth_integrtaion_6_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_29, QB=>nx31350, D=>nx21923, 
      CLK=>clk, R=>rst);
   ix31353 : nand03 port map ( Y=>nx31352, A0=>nx36171, A1=>nx13206, A2=>
      nx35527);
   ix13207 : xnor2 port map ( Y=>nx13206, A0=>nx31355, A1=>nx13312);
   ix31356 : aoi22 port map ( Y=>nx31355, A0=>
      booth_booth_integrtaion_6_booth_output_29, A1=>nx13154, B0=>nx13134, 
      B1=>nx13311);
   ix31359 : nor02ii port map ( Y=>nx31358, A0=>nx13120, A1=>
      mdr_data_out(125));
   ix13121 : nor02ii port map ( Y=>nx13120, A0=>mdr_data_out(124), A1=>
      nx13096);
   ix13145 : nor02ii port map ( Y=>nx13144, A0=>mdr_data_out(125), A1=>
      nx13120);
   ix31369 : xnor2 port map ( Y=>nx31368, A0=>nx13182, A1=>nx13192);
   ix13183 : oai22 port map ( Y=>nx13182, A0=>nx31355, A1=>nx31371, B0=>
      nx31380, B1=>nx35549);
   ix31374 : aoi32 port map ( Y=>nx31373, A0=>nx13164, A1=>nx35027, A2=>
      nx31378, B0=>mdr_data_out(126), B1=>nx35021);
   ix13165 : nand02 port map ( Y=>nx13164, A0=>nx31376, A1=>
      mdr_data_out(126));
   booth_booth_integrtaion_6_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_31, QB=>nx31380, D=>nx21913, 
      CLK=>clk, R=>rst);
   ix31384 : aoi22 port map ( Y=>nx31383, A0=>mdr_data_out(127), A1=>nx35021, 
      B0=>nx35027, B1=>nx13184);
   ix13185 : xnor2 port map ( Y=>nx13184, A0=>mdr_data_out(127), A1=>nx13168
   );
   ix13169 : nor02ii port map ( Y=>nx13168, A0=>mdr_data_out(126), A1=>
      nx13144);
   ix31388 : aoi32 port map ( Y=>nx31387, A0=>nx13140, A1=>nx35027, A2=>
      nx31376, B0=>mdr_data_out(125), B1=>nx35021);
   ix31391 : aoi32 port map ( Y=>nx31390, A0=>nx13092, A1=>nx35027, A2=>
      nx31341, B0=>mdr_data_out(123), B1=>nx35021);
   ix31394 : aoi32 port map ( Y=>nx31393, A0=>nx13044, A1=>nx35027, A2=>
      nx31306, B0=>mdr_data_out(121), B1=>nx35021);
   ix31397 : aoi32 port map ( Y=>nx31396, A0=>nx12996, A1=>nx35027, A2=>
      nx31271, B0=>mdr_data_out(119), B1=>nx35021);
   ix31400 : aoi32 port map ( Y=>nx31399, A0=>nx12948, A1=>nx35027, A2=>
      nx31236, B0=>mdr_data_out(117), B1=>nx35021);
   ix31403 : aoi32 port map ( Y=>nx31402, A0=>nx12900, A1=>nx12836, A2=>
      nx31201, B0=>mdr_data_out(115), B1=>nx35023);
   ix31406 : aoi32 port map ( Y=>nx31405, A0=>nx12850, A1=>nx12836, A2=>
      nx31150, B0=>mdr_data_out(113), B1=>nx35023);
   booth_booth_integrtaion_6_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_6_booth_output_16, QB=>nx31131, D=>nx22053, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_6_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_6_15, QB=>nx31409, D=>nx22063, CLK=>clk, 
      R=>rst);
   ix13575 : aoi21 port map ( Y=>nx13574, A0=>label_7_output(0), A1=>nx35771, 
      B0=>nx35919);
   ix23624 : oai21 port map ( Y=>nx23623, A0=>nx31429, A1=>nx34785, B0=>
      nx31431);
   max_calc_reg_comparator_fourth_inp2_0 : dff port map ( Q=>OPEN, QB=>
      nx31429, D=>nx23623, CLK=>clk);
   ix31432 : nand03 port map ( Y=>nx31431, A0=>label_8_output(0), A1=>
      nx35461, A2=>nx34785);
   labelsregfile_label8_loop1_0_fx_reg_q : dffr port map ( Q=>
      label_8_output(0), QB=>OPEN, D=>nx23073, CLK=>clk, R=>rst);
   lat_label_8_input_0 : latch port map ( Q=>label_8_input_0, D=>nx14902, 
      CLK=>nx34529);
   ix14903 : oai21 port map ( Y=>nx14902, A0=>nx31437, A1=>nx34429, B0=>
      nx31441);
   reg_label_8_input_state_machine_0 : dffr port map ( Q=>
      label_8_input_state_machine_0, QB=>nx31437, D=>nx23063, CLK=>clk, R=>
      rst);
   ix31442 : oai21 port map ( Y=>nx31441, A0=>nx35775, A1=>label_8_output(0), 
      B0=>nx14890);
   booth_booth_integrtaion_7_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_1, QB=>OPEN, D=>nx23043, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_2, QB=>nx31862, D=>nx23033, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_3, QB=>OPEN, D=>nx23023, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_4, QB=>nx31860, D=>nx23013, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_5, QB=>OPEN, D=>nx23003, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_6, QB=>nx31858, D=>nx22993, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_7, QB=>OPEN, D=>nx22983, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_8, QB=>nx31856, D=>nx22973, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_9, QB=>OPEN, D=>nx22963, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_10, QB=>nx31854, D=>nx22953, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_11, QB=>OPEN, D=>nx22943, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_12, QB=>nx31852, D=>nx22933, CLK=>clk, 
      R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_13, QB=>OPEN, D=>nx22923, CLK=>clk, R
      =>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_14, QB=>nx31850, D=>nx22913, CLK=>clk, 
      R=>rst);
   ix31491 : aoi22 port map ( Y=>nx31490, A0=>mdr_data_out(15), A1=>nx35043, 
      B0=>nx14688, B1=>nx14694);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_0_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_reg_output_0, QB=>OPEN, 
      D=>nx22553, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_0, QB=>OPEN, D=>nx22539, CLK
      =>clk, S=>nx34493);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_9_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_reg_output_9, QB=>OPEN, 
      D=>nx22733, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_9, QB=>OPEN, D=>nx22723, CLK
      =>clk, R=>nx34493);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_8_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_8, QB=>OPEN, 
      D=>nx22713, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_8, QB=>OPEN, D=>nx22703, CLK
      =>clk, R=>nx34493);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_7_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_7, QB=>OPEN, 
      D=>nx22693, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_7, QB=>OPEN, D=>nx22683, CLK
      =>clk, R=>nx34493);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_6_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_6, QB=>OPEN, 
      D=>nx22673, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_6, QB=>OPEN, D=>nx22663, CLK
      =>clk, R=>nx34491);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_5_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_5, QB=>OPEN, 
      D=>nx22653, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_5, QB=>OPEN, D=>nx22643, CLK
      =>clk, R=>nx34491);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_4_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_4, QB=>OPEN, 
      D=>nx22633, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_4, QB=>OPEN, D=>nx22623, CLK
      =>clk, R=>nx34491);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_3_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_3, QB=>OPEN, 
      D=>nx22613, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_3, QB=>OPEN, D=>nx22603, CLK
      =>clk, R=>nx34491);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_2_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_2, QB=>OPEN, 
      D=>nx22593, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_2, QB=>OPEN, D=>nx22583, CLK
      =>clk, R=>nx34491);
   booth_booth_integrtaion_7_shift_Reg_Reg_loop1_1_fx_reg_q : dffr
       port map ( Q=>booth_booth_integrtaion_7_shift_Reg_output_1, QB=>OPEN, 
      D=>nx22573, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_booth_integrtaion_7_shift_Reg_count_1, QB=>OPEN, D=>nx22563, CLK
      =>clk, R=>nx34491);
   ix22534 : nand02 port map ( Y=>nx22533, A0=>nx35839, A1=>nx35029);
   booth_booth_integrtaion_7_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, 
      QB=>nx31537, D=>nx22533, CLK=>clk, S=>nx34491);
   ix14689 : nand02 port map ( Y=>nx14688, A0=>nx31558, A1=>nx31570);
   ix31559 : oai21 port map ( Y=>nx31558, A0=>nx35057, A1=>nx35051, B0=>
      mdr_data_out(128));
   ix22744 : oai21 port map ( Y=>nx22743, A0=>nx31563, A1=>nx35551, B0=>
      nx31565);
   booth_booth_integrtaion_7_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx31563, D=>nx22743, CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      OPEN, QB=>nx31567, D=>nx23053, CLK=>clk, R=>rst);
   ix31575 : xnor2 port map ( Y=>nx31574, A0=>nx14158, A1=>nx13334);
   ix22884 : oai21 port map ( Y=>nx22883, A0=>nx31580, A1=>nx35551, B0=>
      nx31582);
   booth_booth_integrtaion_7_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_17, QB=>nx31580, D=>nx22883, 
      CLK=>clk, R=>rst);
   ix31583 : nand03 port map ( Y=>nx31582, A0=>nx35559, A1=>nx14666, A2=>
      nx36179);
   ix14667 : xnor2 port map ( Y=>nx14666, A0=>nx31585, A1=>nx13335);
   ix31586 : aoi22 port map ( Y=>nx31585, A0=>
      booth_booth_integrtaion_7_booth_output_17, A1=>nx14182, B0=>nx14158, 
      B1=>nx13334);
   ix14167 : nand02 port map ( Y=>nx14166, A0=>mdr_data_out(129), A1=>
      mdr_data_out(128));
   ix31590 : or02 port map ( Y=>nx31589, A0=>mdr_data_out(128), A1=>
      mdr_data_out(129));
   ix31596 : xnor2 port map ( Y=>nx31595, A0=>nx14210, A1=>nx13336);
   ix14211 : oai22 port map ( Y=>nx14210, A0=>nx31585, A1=>nx31598, B0=>
      nx31605, B1=>nx35563);
   ix31601 : aoi32 port map ( Y=>nx31600, A0=>nx14192, A1=>nx35057, A2=>
      nx31603, B0=>mdr_data_out(130), B1=>nx35051);
   ix14193 : oai21 port map ( Y=>nx14192, A0=>mdr_data_out(128), A1=>
      mdr_data_out(129), B0=>mdr_data_out(130));
   booth_booth_integrtaion_7_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_18, QB=>nx31605, D=>nx22873, 
      CLK=>clk, R=>rst);
   ix22864 : oai21 port map ( Y=>nx22863, A0=>nx31610, A1=>nx35551, B0=>
      nx31612);
   booth_booth_integrtaion_7_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_19, QB=>nx31610, D=>nx22863, 
      CLK=>clk, R=>rst);
   ix31613 : nand03 port map ( Y=>nx31612, A0=>nx35559, A1=>nx14642, A2=>
      nx36179);
   ix14643 : xnor2 port map ( Y=>nx14642, A0=>nx31615, A1=>nx13337);
   ix31616 : aoi22 port map ( Y=>nx31615, A0=>
      booth_booth_integrtaion_7_booth_output_19, A1=>nx14230, B0=>nx14210, 
      B1=>nx13336);
   ix31619 : nor02ii port map ( Y=>nx31618, A0=>nx14196, A1=>
      mdr_data_out(131));
   ix14197 : nor03_2x port map ( Y=>nx14196, A0=>mdr_data_out(130), A1=>
      mdr_data_out(128), A2=>mdr_data_out(129));
   ix14221 : nor04 port map ( Y=>nx14220, A0=>mdr_data_out(131), A1=>
      mdr_data_out(130), A2=>mdr_data_out(128), A3=>mdr_data_out(129));
   ix31633 : xnor2 port map ( Y=>nx31632, A0=>nx14258, A1=>nx13339);
   ix14259 : oai22 port map ( Y=>nx14258, A0=>nx31615, A1=>nx31635, B0=>
      nx31644, B1=>nx35565);
   ix31638 : aoi32 port map ( Y=>nx31637, A0=>nx14240, A1=>nx35057, A2=>
      nx31642, B0=>mdr_data_out(132), B1=>nx35051);
   ix14241 : nand02 port map ( Y=>nx14240, A0=>nx31640, A1=>
      mdr_data_out(132));
   booth_booth_integrtaion_7_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_20, QB=>nx31644, D=>nx22853, 
      CLK=>clk, R=>rst);
   ix22844 : oai21 port map ( Y=>nx22843, A0=>nx31649, A1=>nx35551, B0=>
      nx31651);
   booth_booth_integrtaion_7_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_21, QB=>nx31649, D=>nx22843, 
      CLK=>clk, R=>rst);
   ix31652 : nand03 port map ( Y=>nx31651, A0=>nx35559, A1=>nx14618, A2=>
      nx36179);
   ix14619 : xnor2 port map ( Y=>nx14618, A0=>nx31654, A1=>nx13341);
   ix31655 : aoi22 port map ( Y=>nx31654, A0=>
      booth_booth_integrtaion_7_booth_output_21, A1=>nx14278, B0=>nx14258, 
      B1=>nx13339);
   ix31658 : nor02ii port map ( Y=>nx31657, A0=>nx14244, A1=>
      mdr_data_out(133));
   ix14245 : nor02ii port map ( Y=>nx14244, A0=>mdr_data_out(132), A1=>
      nx14220);
   ix14269 : nor02ii port map ( Y=>nx14268, A0=>mdr_data_out(133), A1=>
      nx14244);
   ix31668 : xnor2 port map ( Y=>nx31667, A0=>nx14306, A1=>nx13343);
   ix14307 : oai22 port map ( Y=>nx14306, A0=>nx31654, A1=>nx31670, B0=>
      nx31679, B1=>nx35567);
   ix31673 : aoi32 port map ( Y=>nx31672, A0=>nx14288, A1=>nx35057, A2=>
      nx31677, B0=>mdr_data_out(134), B1=>nx35051);
   ix14289 : nand02 port map ( Y=>nx14288, A0=>nx31675, A1=>
      mdr_data_out(134));
   booth_booth_integrtaion_7_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_22, QB=>nx31679, D=>nx22833, 
      CLK=>clk, R=>rst);
   ix22824 : oai21 port map ( Y=>nx22823, A0=>nx31684, A1=>nx35551, B0=>
      nx31686);
   booth_booth_integrtaion_7_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_23, QB=>nx31684, D=>nx22823, 
      CLK=>clk, R=>rst);
   ix31687 : nand03 port map ( Y=>nx31686, A0=>nx35559, A1=>nx14594, A2=>
      nx35553);
   ix14595 : xnor2 port map ( Y=>nx14594, A0=>nx31689, A1=>nx13344);
   ix31690 : aoi22 port map ( Y=>nx31689, A0=>
      booth_booth_integrtaion_7_booth_output_23, A1=>nx14326, B0=>nx14306, 
      B1=>nx13343);
   ix31693 : nor02ii port map ( Y=>nx31692, A0=>nx14292, A1=>
      mdr_data_out(135));
   ix14293 : nor02ii port map ( Y=>nx14292, A0=>mdr_data_out(134), A1=>
      nx14268);
   ix14317 : nor02ii port map ( Y=>nx14316, A0=>mdr_data_out(135), A1=>
      nx14292);
   ix31703 : xnor2 port map ( Y=>nx31702, A0=>nx14354, A1=>nx13345);
   ix14355 : oai22 port map ( Y=>nx14354, A0=>nx31689, A1=>nx31705, B0=>
      nx31714, B1=>nx35569);
   ix31708 : aoi32 port map ( Y=>nx31707, A0=>nx14336, A1=>nx35057, A2=>
      nx31712, B0=>mdr_data_out(136), B1=>nx35051);
   ix14337 : nand02 port map ( Y=>nx14336, A0=>nx31710, A1=>
      mdr_data_out(136));
   booth_booth_integrtaion_7_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_24, QB=>nx31714, D=>nx22813, 
      CLK=>clk, R=>rst);
   ix22804 : oai21 port map ( Y=>nx22803, A0=>nx31719, A1=>nx35553, B0=>
      nx31721);
   booth_booth_integrtaion_7_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_25, QB=>nx31719, D=>nx22803, 
      CLK=>clk, R=>rst);
   ix31722 : nand03 port map ( Y=>nx31721, A0=>nx35559, A1=>nx14570, A2=>
      nx35553);
   ix14571 : xnor2 port map ( Y=>nx14570, A0=>nx31724, A1=>nx13346);
   ix31725 : aoi22 port map ( Y=>nx31724, A0=>
      booth_booth_integrtaion_7_booth_output_25, A1=>nx14374, B0=>nx14354, 
      B1=>nx13345);
   ix31728 : nor02ii port map ( Y=>nx31727, A0=>nx14340, A1=>
      mdr_data_out(137));
   ix14341 : nor02ii port map ( Y=>nx14340, A0=>mdr_data_out(136), A1=>
      nx14316);
   ix14365 : nor02ii port map ( Y=>nx14364, A0=>mdr_data_out(137), A1=>
      nx14340);
   ix31738 : xnor2 port map ( Y=>nx31737, A0=>nx14402, A1=>nx13347);
   ix14403 : oai22 port map ( Y=>nx14402, A0=>nx31724, A1=>nx31740, B0=>
      nx31749, B1=>nx35571);
   ix31743 : aoi32 port map ( Y=>nx31742, A0=>nx14384, A1=>nx35057, A2=>
      nx31747, B0=>mdr_data_out(138), B1=>nx35051);
   ix14385 : nand02 port map ( Y=>nx14384, A0=>nx31745, A1=>
      mdr_data_out(138));
   booth_booth_integrtaion_7_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_26, QB=>nx31749, D=>nx22793, 
      CLK=>clk, R=>rst);
   ix22784 : oai21 port map ( Y=>nx22783, A0=>nx31754, A1=>nx35553, B0=>
      nx31756);
   booth_booth_integrtaion_7_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_27, QB=>nx31754, D=>nx22783, 
      CLK=>clk, R=>rst);
   ix31757 : nand03 port map ( Y=>nx31756, A0=>nx35559, A1=>nx14546, A2=>
      nx35553);
   ix14547 : xnor2 port map ( Y=>nx14546, A0=>nx31759, A1=>nx13348);
   ix31760 : aoi22 port map ( Y=>nx31759, A0=>
      booth_booth_integrtaion_7_booth_output_27, A1=>nx14422, B0=>nx14402, 
      B1=>nx13347);
   ix31763 : nor02ii port map ( Y=>nx31762, A0=>nx14388, A1=>
      mdr_data_out(139));
   ix14389 : nor02ii port map ( Y=>nx14388, A0=>mdr_data_out(138), A1=>
      nx14364);
   ix14413 : nor02ii port map ( Y=>nx14412, A0=>mdr_data_out(139), A1=>
      nx14388);
   ix31773 : xnor2 port map ( Y=>nx31772, A0=>nx14450, A1=>nx13349);
   ix14451 : oai22 port map ( Y=>nx14450, A0=>nx31759, A1=>nx31775, B0=>
      nx31784, B1=>nx35573);
   ix31778 : aoi32 port map ( Y=>nx31777, A0=>nx14432, A1=>nx35057, A2=>
      nx31782, B0=>mdr_data_out(140), B1=>nx35051);
   ix14433 : nand02 port map ( Y=>nx14432, A0=>nx31780, A1=>
      mdr_data_out(140));
   booth_booth_integrtaion_7_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_28, QB=>nx31784, D=>nx22773, 
      CLK=>clk, R=>rst);
   ix22764 : oai21 port map ( Y=>nx22763, A0=>nx31789, A1=>nx35553, B0=>
      nx31791);
   booth_booth_integrtaion_7_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_29, QB=>nx31789, D=>nx22763, 
      CLK=>clk, R=>rst);
   ix31792 : nand03 port map ( Y=>nx31791, A0=>nx36187, A1=>nx14522, A2=>
      nx35553);
   ix14523 : xnor2 port map ( Y=>nx14522, A0=>nx31794, A1=>nx13351);
   ix31795 : aoi22 port map ( Y=>nx31794, A0=>
      booth_booth_integrtaion_7_booth_output_29, A1=>nx14470, B0=>nx14450, 
      B1=>nx13349);
   ix31798 : nor02ii port map ( Y=>nx31797, A0=>nx14436, A1=>
      mdr_data_out(141));
   ix14437 : nor02ii port map ( Y=>nx14436, A0=>mdr_data_out(140), A1=>
      nx14412);
   ix14461 : nor02ii port map ( Y=>nx14460, A0=>mdr_data_out(141), A1=>
      nx14436);
   ix31808 : xnor2 port map ( Y=>nx31807, A0=>nx14498, A1=>nx14508);
   ix14499 : oai22 port map ( Y=>nx14498, A0=>nx31794, A1=>nx31810, B0=>
      nx31819, B1=>nx35575);
   ix31813 : aoi32 port map ( Y=>nx31812, A0=>nx14480, A1=>nx35059, A2=>
      nx31817, B0=>mdr_data_out(142), B1=>nx35053);
   ix14481 : nand02 port map ( Y=>nx14480, A0=>nx31815, A1=>
      mdr_data_out(142));
   booth_booth_integrtaion_7_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_31, QB=>nx31819, D=>nx22753, 
      CLK=>clk, R=>rst);
   ix31823 : aoi22 port map ( Y=>nx31822, A0=>mdr_data_out(143), A1=>nx35053, 
      B0=>nx35059, B1=>nx14500);
   ix14501 : xnor2 port map ( Y=>nx14500, A0=>mdr_data_out(143), A1=>nx14484
   );
   ix14485 : nor02ii port map ( Y=>nx14484, A0=>mdr_data_out(142), A1=>
      nx14460);
   ix31827 : aoi32 port map ( Y=>nx31826, A0=>nx14456, A1=>nx35059, A2=>
      nx31815, B0=>mdr_data_out(141), B1=>nx35053);
   ix31830 : aoi32 port map ( Y=>nx31829, A0=>nx14408, A1=>nx35059, A2=>
      nx31780, B0=>mdr_data_out(139), B1=>nx35053);
   ix31833 : aoi32 port map ( Y=>nx31832, A0=>nx14360, A1=>nx35059, A2=>
      nx31745, B0=>mdr_data_out(137), B1=>nx35053);
   ix31836 : aoi32 port map ( Y=>nx31835, A0=>nx14312, A1=>nx35059, A2=>
      nx31710, B0=>mdr_data_out(135), B1=>nx35053);
   ix31839 : aoi32 port map ( Y=>nx31838, A0=>nx14264, A1=>nx35059, A2=>
      nx31675, B0=>mdr_data_out(133), B1=>nx35053);
   ix31842 : aoi32 port map ( Y=>nx31841, A0=>nx14216, A1=>nx14152, A2=>
      nx31640, B0=>mdr_data_out(131), B1=>nx35055);
   ix31845 : aoi32 port map ( Y=>nx31844, A0=>nx14166, A1=>nx14152, A2=>
      nx31589, B0=>mdr_data_out(129), B1=>nx35055);
   booth_booth_integrtaion_7_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_booth_integrtaion_7_booth_output_16, QB=>nx31570, D=>nx22893, 
      CLK=>clk, R=>rst);
   booth_booth_integrtaion_7_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_booth_integration_output_7_15, QB=>nx31848, D=>nx22903, CLK=>clk, 
      R=>rst);
   ix14891 : aoi21 port map ( Y=>nx14890, A0=>label_8_output(0), A1=>nx35775, 
      B0=>nx35919);
   ix15875 : xnor2 port map ( Y=>nx15874, A0=>nx31867, A1=>nx15872);
   ix31868 : aoi22 port map ( Y=>nx31867, A0=>nx31869, A1=>
      max_calc_comparator_fourth_inp1_14, B0=>nx15360, B1=>nx15778);
   max_calc_reg_comparator_fourth_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx31869, D=>nx23353, CLK=>clk);
   ix23354 : oai21 port map ( Y=>nx23353, A0=>nx31869, A1=>nx34785, B0=>
      nx31872);
   labelsregfile_label8_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_8_output(14), QB=>nx32056, D=>nx23343, CLK=>clk, R=>rst);
   lat_label_8_input_14 : latch port map ( Q=>label_8_input_14, D=>nx15338, 
      CLK=>nx34533);
   reg_label_8_input_state_machine_14 : dffr port map ( Q=>
      label_8_input_state_machine_14, QB=>OPEN, D=>nx22523, CLK=>clk, R=>rst
   );
   ix15335 : xor2 port map ( Y=>nx15334, A0=>nx31882, A1=>nx32054);
   ix31883 : aoi22 port map ( Y=>nx31882, A0=>label_8_output(13), A1=>
      booth_booth_integration_output_7_13, B0=>nx15298, B1=>nx13370);
   labelsregfile_label8_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_8_output(13), QB=>OPEN, D=>nx23333, CLK=>clk, R=>rst);
   lat_label_8_input_13 : latch port map ( Q=>label_8_input_13, D=>nx15312, 
      CLK=>nx34533);
   reg_label_8_input_state_machine_13 : dffr port map ( Q=>
      label_8_input_state_machine_13, QB=>OPEN, D=>nx23323, CLK=>clk, R=>rst
   );
   ix15309 : xnor2 port map ( Y=>nx15308, A0=>nx15298, A1=>nx32050);
   ix15299 : oai22 port map ( Y=>nx15298, A0=>nx31893, A1=>nx32039, B0=>
      nx32049, B1=>nx31852);
   ix31894 : aoi22 port map ( Y=>nx31893, A0=>label_8_output(11), A1=>
      booth_booth_integration_output_7_11, B0=>nx15234, B1=>nx13368);
   labelsregfile_label8_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_8_output(11), QB=>OPEN, D=>nx23293, CLK=>clk, R=>rst);
   lat_label_8_input_11 : latch port map ( Q=>label_8_input_11, D=>nx15248, 
      CLK=>nx34533);
   reg_label_8_input_state_machine_11 : dffr port map ( Q=>
      label_8_input_state_machine_11, QB=>OPEN, D=>nx23283, CLK=>clk, R=>rst
   );
   ix15245 : xnor2 port map ( Y=>nx15244, A0=>nx15234, A1=>nx32035);
   ix15235 : oai22 port map ( Y=>nx15234, A0=>nx31904, A1=>nx32024, B0=>
      nx32034, B1=>nx31854);
   ix31905 : aoi22 port map ( Y=>nx31904, A0=>label_8_output(9), A1=>
      booth_booth_integration_output_7_9, B0=>nx15170, B1=>nx13365);
   labelsregfile_label8_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_8_output(9), QB=>OPEN, D=>nx23253, CLK=>clk, R=>rst);
   lat_label_8_input_9 : latch port map ( Q=>label_8_input_9, D=>nx15184, 
      CLK=>nx34533);
   reg_label_8_input_state_machine_9 : dffr port map ( Q=>
      label_8_input_state_machine_9, QB=>OPEN, D=>nx23243, CLK=>clk, R=>rst
   );
   ix15181 : xnor2 port map ( Y=>nx15180, A0=>nx15170, A1=>nx32020);
   ix15171 : oai22 port map ( Y=>nx15170, A0=>nx31915, A1=>nx32009, B0=>
      nx32019, B1=>nx31856);
   ix31916 : aoi22 port map ( Y=>nx31915, A0=>label_8_output(7), A1=>
      booth_booth_integration_output_7_7, B0=>nx15106, B1=>nx13361);
   labelsregfile_label8_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_8_output(7), QB=>OPEN, D=>nx23213, CLK=>clk, R=>rst);
   lat_label_8_input_7 : latch port map ( Q=>label_8_input_7, D=>nx15120, 
      CLK=>nx34531);
   reg_label_8_input_state_machine_7 : dffr port map ( Q=>
      label_8_input_state_machine_7, QB=>OPEN, D=>nx23203, CLK=>clk, R=>rst
   );
   ix15117 : xnor2 port map ( Y=>nx15116, A0=>nx15106, A1=>nx32005);
   ix15107 : oai22 port map ( Y=>nx15106, A0=>nx31926, A1=>nx31994, B0=>
      nx32004, B1=>nx31858);
   ix31927 : aoi22 port map ( Y=>nx31926, A0=>label_8_output(5), A1=>
      booth_booth_integration_output_7_5, B0=>nx15042, B1=>nx13359);
   labelsregfile_label8_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_8_output(5), QB=>OPEN, D=>nx23173, CLK=>clk, R=>rst);
   lat_label_8_input_5 : latch port map ( Q=>label_8_input_5, D=>nx15056, 
      CLK=>nx34531);
   reg_label_8_input_state_machine_5 : dffr port map ( Q=>
      label_8_input_state_machine_5, QB=>OPEN, D=>nx23163, CLK=>clk, R=>rst
   );
   ix15053 : xnor2 port map ( Y=>nx15052, A0=>nx15042, A1=>nx31990);
   ix15043 : oai22 port map ( Y=>nx15042, A0=>nx31937, A1=>nx31979, B0=>
      nx31989, B1=>nx31860);
   ix31938 : aoi22 port map ( Y=>nx31937, A0=>label_8_output(3), A1=>
      booth_booth_integration_output_7_3, B0=>nx14978, B1=>nx13357);
   labelsregfile_label8_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_8_output(3), QB=>OPEN, D=>nx23133, CLK=>clk, R=>rst);
   lat_label_8_input_3 : latch port map ( Q=>label_8_input_3, D=>nx14992, 
      CLK=>nx34531);
   reg_label_8_input_state_machine_3 : dffr port map ( Q=>
      label_8_input_state_machine_3, QB=>OPEN, D=>nx23123, CLK=>clk, R=>rst
   );
   ix14989 : xnor2 port map ( Y=>nx14988, A0=>nx14978, A1=>nx31975);
   ix14979 : oai22 port map ( Y=>nx14978, A0=>nx31948, A1=>nx31964, B0=>
      nx31974, B1=>nx31862);
   ix31949 : aoi32 port map ( Y=>nx31948, A0=>label_8_output(0), A1=>nx35775, 
      A2=>nx13355, B0=>label_8_output(1), B1=>
      booth_booth_integration_output_7_1);
   labelsregfile_label8_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_8_output(1), QB=>OPEN, D=>nx23093, CLK=>clk, R=>rst);
   lat_label_8_input_1 : latch port map ( Q=>label_8_input_1, D=>nx14928, 
      CLK=>nx34531);
   reg_label_8_input_state_machine_1 : dffr port map ( Q=>
      label_8_input_state_machine_1, QB=>OPEN, D=>nx23083, CLK=>clk, R=>rst
   );
   ix14925 : xor2 port map ( Y=>nx14924, A0=>nx31959, A1=>nx31961);
   ix31960 : nand02 port map ( Y=>nx31959, A0=>label_8_output(0), A1=>
      nx35775);
   ix31962 : xnor2 port map ( Y=>nx31961, A0=>
      booth_booth_integration_output_7_1, A1=>label_8_output(1));
   labelsregfile_label8_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_8_output(2), QB=>nx31974, D=>nx23113, CLK=>clk, R=>rst);
   lat_label_8_input_2 : latch port map ( Q=>label_8_input_2, D=>nx14960, 
      CLK=>nx34531);
   reg_label_8_input_state_machine_2 : dffr port map ( Q=>
      label_8_input_state_machine_2, QB=>OPEN, D=>nx23103, CLK=>clk, R=>rst
   );
   ix14957 : xor2 port map ( Y=>nx14956, A0=>nx31948, A1=>nx31964);
   ix31976 : xnor2 port map ( Y=>nx31975, A0=>
      booth_booth_integration_output_7_3, A1=>label_8_output(3));
   labelsregfile_label8_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_8_output(4), QB=>nx31989, D=>nx23153, CLK=>clk, R=>rst);
   lat_label_8_input_4 : latch port map ( Q=>label_8_input_4, D=>nx15024, 
      CLK=>nx34531);
   reg_label_8_input_state_machine_4 : dffr port map ( Q=>
      label_8_input_state_machine_4, QB=>OPEN, D=>nx23143, CLK=>clk, R=>rst
   );
   ix15021 : xor2 port map ( Y=>nx15020, A0=>nx31937, A1=>nx31979);
   ix31991 : xnor2 port map ( Y=>nx31990, A0=>
      booth_booth_integration_output_7_5, A1=>label_8_output(5));
   labelsregfile_label8_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_8_output(6), QB=>nx32004, D=>nx23193, CLK=>clk, R=>rst);
   lat_label_8_input_6 : latch port map ( Q=>label_8_input_6, D=>nx15088, 
      CLK=>nx34531);
   reg_label_8_input_state_machine_6 : dffr port map ( Q=>
      label_8_input_state_machine_6, QB=>OPEN, D=>nx23183, CLK=>clk, R=>rst
   );
   ix15085 : xor2 port map ( Y=>nx15084, A0=>nx31926, A1=>nx31994);
   ix32006 : xnor2 port map ( Y=>nx32005, A0=>
      booth_booth_integration_output_7_7, A1=>label_8_output(7));
   labelsregfile_label8_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_8_output(8), QB=>nx32019, D=>nx23233, CLK=>clk, R=>rst);
   lat_label_8_input_8 : latch port map ( Q=>label_8_input_8, D=>nx15152, 
      CLK=>nx34533);
   reg_label_8_input_state_machine_8 : dffr port map ( Q=>
      label_8_input_state_machine_8, QB=>OPEN, D=>nx23223, CLK=>clk, R=>rst
   );
   ix15149 : xor2 port map ( Y=>nx15148, A0=>nx31915, A1=>nx32009);
   ix32021 : xnor2 port map ( Y=>nx32020, A0=>
      booth_booth_integration_output_7_9, A1=>label_8_output(9));
   labelsregfile_label8_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_8_output(10), QB=>nx32034, D=>nx23273, CLK=>clk, R=>rst);
   lat_label_8_input_10 : latch port map ( Q=>label_8_input_10, D=>nx15216, 
      CLK=>nx34533);
   reg_label_8_input_state_machine_10 : dffr port map ( Q=>
      label_8_input_state_machine_10, QB=>OPEN, D=>nx23263, CLK=>clk, R=>rst
   );
   ix15213 : xor2 port map ( Y=>nx15212, A0=>nx31904, A1=>nx32024);
   ix32036 : xnor2 port map ( Y=>nx32035, A0=>
      booth_booth_integration_output_7_11, A1=>label_8_output(11));
   labelsregfile_label8_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_8_output(12), QB=>nx32049, D=>nx23313, CLK=>clk, R=>rst);
   lat_label_8_input_12 : latch port map ( Q=>label_8_input_12, D=>nx15280, 
      CLK=>nx34533);
   reg_label_8_input_state_machine_12 : dffr port map ( Q=>
      label_8_input_state_machine_12, QB=>OPEN, D=>nx23303, CLK=>clk, R=>rst
   );
   ix15277 : xor2 port map ( Y=>nx15276, A0=>nx31893, A1=>nx32039);
   ix32051 : xnor2 port map ( Y=>nx32050, A0=>
      booth_booth_integration_output_7_13, A1=>label_8_output(13));
   ix22514 : oai21 port map ( Y=>nx22513, A0=>nx32059, A1=>nx34785, B0=>
      nx32061);
   max_calc_reg_comparator_fourth_inp1_14 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_14, QB=>nx32059, D=>nx22513, CLK=>clk
   );
   labelsregfile_label7_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_7_output(14), QB=>nx32245, D=>nx22503, CLK=>clk, R=>rst);
   lat_label_7_input_14 : latch port map ( Q=>label_7_input_14, D=>nx14022, 
      CLK=>nx34537);
   reg_label_7_input_state_machine_14 : dffr port map ( Q=>
      label_7_input_state_machine_14, QB=>OPEN, D=>nx21683, CLK=>clk, R=>rst
   );
   ix14019 : xor2 port map ( Y=>nx14018, A0=>nx32071, A1=>nx32243);
   ix32072 : aoi22 port map ( Y=>nx32071, A0=>label_7_output(13), A1=>
      booth_booth_integration_output_6_13, B0=>nx13982, B1=>nx13332);
   labelsregfile_label7_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_7_output(13), QB=>OPEN, D=>nx22493, CLK=>clk, R=>rst);
   lat_label_7_input_13 : latch port map ( Q=>label_7_input_13, D=>nx13996, 
      CLK=>nx34537);
   reg_label_7_input_state_machine_13 : dffr port map ( Q=>
      label_7_input_state_machine_13, QB=>OPEN, D=>nx22483, CLK=>clk, R=>rst
   );
   ix13993 : xnor2 port map ( Y=>nx13992, A0=>nx13982, A1=>nx32239);
   ix13983 : oai22 port map ( Y=>nx13982, A0=>nx32082, A1=>nx32228, B0=>
      nx32238, B1=>nx31413);
   ix32083 : aoi22 port map ( Y=>nx32082, A0=>label_7_output(11), A1=>
      booth_booth_integration_output_6_11, B0=>nx13918, B1=>nx13329);
   labelsregfile_label7_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_7_output(11), QB=>OPEN, D=>nx22453, CLK=>clk, R=>rst);
   lat_label_7_input_11 : latch port map ( Q=>label_7_input_11, D=>nx13932, 
      CLK=>nx34537);
   reg_label_7_input_state_machine_11 : dffr port map ( Q=>
      label_7_input_state_machine_11, QB=>OPEN, D=>nx22443, CLK=>clk, R=>rst
   );
   ix13929 : xnor2 port map ( Y=>nx13928, A0=>nx13918, A1=>nx32224);
   ix13919 : oai22 port map ( Y=>nx13918, A0=>nx32093, A1=>nx32213, B0=>
      nx32223, B1=>nx31415);
   ix32094 : aoi22 port map ( Y=>nx32093, A0=>label_7_output(9), A1=>
      booth_booth_integration_output_6_9, B0=>nx13854, B1=>nx13325);
   labelsregfile_label7_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_7_output(9), QB=>OPEN, D=>nx22413, CLK=>clk, R=>rst);
   lat_label_7_input_9 : latch port map ( Q=>label_7_input_9, D=>nx13868, 
      CLK=>nx34537);
   reg_label_7_input_state_machine_9 : dffr port map ( Q=>
      label_7_input_state_machine_9, QB=>OPEN, D=>nx22403, CLK=>clk, R=>rst
   );
   ix13865 : xnor2 port map ( Y=>nx13864, A0=>nx13854, A1=>nx32209);
   ix13855 : oai22 port map ( Y=>nx13854, A0=>nx32104, A1=>nx32198, B0=>
      nx32208, B1=>nx31417);
   ix32105 : aoi22 port map ( Y=>nx32104, A0=>label_7_output(7), A1=>
      booth_booth_integration_output_6_7, B0=>nx13790, B1=>nx13323);
   labelsregfile_label7_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_7_output(7), QB=>OPEN, D=>nx22373, CLK=>clk, R=>rst);
   lat_label_7_input_7 : latch port map ( Q=>label_7_input_7, D=>nx13804, 
      CLK=>nx34535);
   reg_label_7_input_state_machine_7 : dffr port map ( Q=>
      label_7_input_state_machine_7, QB=>OPEN, D=>nx22363, CLK=>clk, R=>rst
   );
   ix13801 : xnor2 port map ( Y=>nx13800, A0=>nx13790, A1=>nx32194);
   ix13791 : oai22 port map ( Y=>nx13790, A0=>nx32115, A1=>nx32183, B0=>
      nx32193, B1=>nx31419);
   ix32116 : aoi22 port map ( Y=>nx32115, A0=>label_7_output(5), A1=>
      booth_booth_integration_output_6_5, B0=>nx13726, B1=>nx13321);
   labelsregfile_label7_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_7_output(5), QB=>OPEN, D=>nx22333, CLK=>clk, R=>rst);
   lat_label_7_input_5 : latch port map ( Q=>label_7_input_5, D=>nx13740, 
      CLK=>nx34535);
   reg_label_7_input_state_machine_5 : dffr port map ( Q=>
      label_7_input_state_machine_5, QB=>OPEN, D=>nx22323, CLK=>clk, R=>rst
   );
   ix13737 : xnor2 port map ( Y=>nx13736, A0=>nx13726, A1=>nx32179);
   ix13727 : oai22 port map ( Y=>nx13726, A0=>nx32126, A1=>nx32168, B0=>
      nx32178, B1=>nx31421);
   ix32127 : aoi22 port map ( Y=>nx32126, A0=>label_7_output(3), A1=>
      booth_booth_integration_output_6_3, B0=>nx13662, B1=>nx13319);
   labelsregfile_label7_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_7_output(3), QB=>OPEN, D=>nx22293, CLK=>clk, R=>rst);
   lat_label_7_input_3 : latch port map ( Q=>label_7_input_3, D=>nx13676, 
      CLK=>nx34535);
   reg_label_7_input_state_machine_3 : dffr port map ( Q=>
      label_7_input_state_machine_3, QB=>OPEN, D=>nx22283, CLK=>clk, R=>rst
   );
   ix13673 : xnor2 port map ( Y=>nx13672, A0=>nx13662, A1=>nx32164);
   ix13663 : oai22 port map ( Y=>nx13662, A0=>nx32137, A1=>nx32153, B0=>
      nx32163, B1=>nx31423);
   ix32138 : aoi32 port map ( Y=>nx32137, A0=>label_7_output(0), A1=>nx35771, 
      A2=>nx13315, B0=>label_7_output(1), B1=>
      booth_booth_integration_output_6_1);
   labelsregfile_label7_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_7_output(1), QB=>OPEN, D=>nx22253, CLK=>clk, R=>rst);
   lat_label_7_input_1 : latch port map ( Q=>label_7_input_1, D=>nx13612, 
      CLK=>nx34535);
   reg_label_7_input_state_machine_1 : dffr port map ( Q=>
      label_7_input_state_machine_1, QB=>OPEN, D=>nx22243, CLK=>clk, R=>rst
   );
   ix13609 : xor2 port map ( Y=>nx13608, A0=>nx32148, A1=>nx32150);
   ix32149 : nand02 port map ( Y=>nx32148, A0=>label_7_output(0), A1=>
      nx35771);
   ix32151 : xnor2 port map ( Y=>nx32150, A0=>
      booth_booth_integration_output_6_1, A1=>label_7_output(1));
   labelsregfile_label7_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_7_output(2), QB=>nx32163, D=>nx22273, CLK=>clk, R=>rst);
   lat_label_7_input_2 : latch port map ( Q=>label_7_input_2, D=>nx13644, 
      CLK=>nx34535);
   reg_label_7_input_state_machine_2 : dffr port map ( Q=>
      label_7_input_state_machine_2, QB=>OPEN, D=>nx22263, CLK=>clk, R=>rst
   );
   ix13641 : xor2 port map ( Y=>nx13640, A0=>nx32137, A1=>nx32153);
   ix32165 : xnor2 port map ( Y=>nx32164, A0=>
      booth_booth_integration_output_6_3, A1=>label_7_output(3));
   labelsregfile_label7_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_7_output(4), QB=>nx32178, D=>nx22313, CLK=>clk, R=>rst);
   lat_label_7_input_4 : latch port map ( Q=>label_7_input_4, D=>nx13708, 
      CLK=>nx34535);
   reg_label_7_input_state_machine_4 : dffr port map ( Q=>
      label_7_input_state_machine_4, QB=>OPEN, D=>nx22303, CLK=>clk, R=>rst
   );
   ix13705 : xor2 port map ( Y=>nx13704, A0=>nx32126, A1=>nx32168);
   ix32180 : xnor2 port map ( Y=>nx32179, A0=>
      booth_booth_integration_output_6_5, A1=>label_7_output(5));
   labelsregfile_label7_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_7_output(6), QB=>nx32193, D=>nx22353, CLK=>clk, R=>rst);
   lat_label_7_input_6 : latch port map ( Q=>label_7_input_6, D=>nx13772, 
      CLK=>nx34535);
   reg_label_7_input_state_machine_6 : dffr port map ( Q=>
      label_7_input_state_machine_6, QB=>OPEN, D=>nx22343, CLK=>clk, R=>rst
   );
   ix13769 : xor2 port map ( Y=>nx13768, A0=>nx32115, A1=>nx32183);
   ix32195 : xnor2 port map ( Y=>nx32194, A0=>
      booth_booth_integration_output_6_7, A1=>label_7_output(7));
   labelsregfile_label7_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_7_output(8), QB=>nx32208, D=>nx22393, CLK=>clk, R=>rst);
   lat_label_7_input_8 : latch port map ( Q=>label_7_input_8, D=>nx13836, 
      CLK=>nx34537);
   reg_label_7_input_state_machine_8 : dffr port map ( Q=>
      label_7_input_state_machine_8, QB=>OPEN, D=>nx22383, CLK=>clk, R=>rst
   );
   ix13833 : xor2 port map ( Y=>nx13832, A0=>nx32104, A1=>nx32198);
   ix32210 : xnor2 port map ( Y=>nx32209, A0=>
      booth_booth_integration_output_6_9, A1=>label_7_output(9));
   labelsregfile_label7_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_7_output(10), QB=>nx32223, D=>nx22433, CLK=>clk, R=>rst);
   lat_label_7_input_10 : latch port map ( Q=>label_7_input_10, D=>nx13900, 
      CLK=>nx34537);
   reg_label_7_input_state_machine_10 : dffr port map ( Q=>
      label_7_input_state_machine_10, QB=>OPEN, D=>nx22423, CLK=>clk, R=>rst
   );
   ix13897 : xor2 port map ( Y=>nx13896, A0=>nx32093, A1=>nx32213);
   ix32225 : xnor2 port map ( Y=>nx32224, A0=>
      booth_booth_integration_output_6_11, A1=>label_7_output(11));
   labelsregfile_label7_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_7_output(12), QB=>nx32238, D=>nx22473, CLK=>clk, R=>rst);
   lat_label_7_input_12 : latch port map ( Q=>label_7_input_12, D=>nx13964, 
      CLK=>nx34537);
   reg_label_7_input_state_machine_12 : dffr port map ( Q=>
      label_7_input_state_machine_12, QB=>OPEN, D=>nx22463, CLK=>clk, R=>rst
   );
   ix13961 : xor2 port map ( Y=>nx13960, A0=>nx32082, A1=>nx32228);
   ix32240 : xnor2 port map ( Y=>nx32239, A0=>
      booth_booth_integration_output_6_13, A1=>label_7_output(13));
   ix15779 : oai22 port map ( Y=>nx15778, A0=>nx32248, A1=>nx32261, B0=>
      max_calc_comparator_fourth_inp2_13, B1=>nx32256);
   ix23364 : oai21 port map ( Y=>nx23363, A0=>nx32252, A1=>nx34785, B0=>
      nx32254);
   max_calc_reg_comparator_fourth_inp2_13 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_13, QB=>nx32252, D=>nx23363, CLK=>clk
   );
   ix32255 : nand03 port map ( Y=>nx32254, A0=>label_8_output(13), A1=>
      nx35463, A2=>nx34787);
   max_calc_reg_comparator_fourth_inp1_13 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_13, QB=>nx32256, D=>nx23373, CLK=>clk
   );
   ix23374 : oai21 port map ( Y=>nx23373, A0=>nx32256, A1=>nx34787, B0=>
      nx32259);
   ix32260 : nand03 port map ( Y=>nx32259, A0=>label_7_output(13), A1=>
      nx35463, A2=>nx34787);
   ix32262 : aoi22 port map ( Y=>nx32261, A0=>nx32263, A1=>
      max_calc_comparator_fourth_inp1_12, B0=>nx15404, B1=>nx15762);
   max_calc_reg_comparator_fourth_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx32263, D=>nx23383, CLK=>clk);
   ix23384 : oai21 port map ( Y=>nx23383, A0=>nx32263, A1=>nx34787, B0=>
      nx32266);
   ix23394 : oai21 port map ( Y=>nx23393, A0=>nx32270, A1=>nx34787, B0=>
      nx32272);
   max_calc_reg_comparator_fourth_inp1_12 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_12, QB=>nx32270, D=>nx23393, CLK=>clk
   );
   ix15763 : oai22 port map ( Y=>nx15762, A0=>nx32276, A1=>nx32289, B0=>
      max_calc_comparator_fourth_inp2_11, B1=>nx32284);
   ix23404 : oai21 port map ( Y=>nx23403, A0=>nx32280, A1=>nx34789, B0=>
      nx32282);
   max_calc_reg_comparator_fourth_inp2_11 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_11, QB=>nx32280, D=>nx23403, CLK=>clk
   );
   ix32283 : nand03 port map ( Y=>nx32282, A0=>label_8_output(11), A1=>
      nx35463, A2=>nx34789);
   max_calc_reg_comparator_fourth_inp1_11 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_11, QB=>nx32284, D=>nx23413, CLK=>clk
   );
   ix23414 : oai21 port map ( Y=>nx23413, A0=>nx32284, A1=>nx34789, B0=>
      nx32287);
   ix32288 : nand03 port map ( Y=>nx32287, A0=>label_7_output(11), A1=>
      nx35463, A2=>nx34789);
   ix32290 : aoi22 port map ( Y=>nx32289, A0=>nx32291, A1=>
      max_calc_comparator_fourth_inp1_10, B0=>nx15448, B1=>nx15746);
   max_calc_reg_comparator_fourth_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx32291, D=>nx23423, CLK=>clk);
   ix23424 : oai21 port map ( Y=>nx23423, A0=>nx32291, A1=>nx34789, B0=>
      nx32294);
   ix23434 : oai21 port map ( Y=>nx23433, A0=>nx32298, A1=>nx34789, B0=>
      nx32300);
   max_calc_reg_comparator_fourth_inp1_10 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_10, QB=>nx32298, D=>nx23433, CLK=>clk
   );
   ix15747 : oai22 port map ( Y=>nx15746, A0=>nx32304, A1=>nx32317, B0=>
      max_calc_comparator_fourth_inp2_9, B1=>nx32312);
   ix23444 : oai21 port map ( Y=>nx23443, A0=>nx32308, A1=>nx34791, B0=>
      nx32310);
   max_calc_reg_comparator_fourth_inp2_9 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_9, QB=>nx32308, D=>nx23443, CLK=>clk);
   ix32311 : nand03 port map ( Y=>nx32310, A0=>label_8_output(9), A1=>
      nx35465, A2=>nx34791);
   max_calc_reg_comparator_fourth_inp1_9 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_9, QB=>nx32312, D=>nx23453, CLK=>clk);
   ix23454 : oai21 port map ( Y=>nx23453, A0=>nx32312, A1=>nx34791, B0=>
      nx32315);
   ix32316 : nand03 port map ( Y=>nx32315, A0=>label_7_output(9), A1=>
      nx35465, A2=>nx34791);
   ix32318 : aoi22 port map ( Y=>nx32317, A0=>nx32319, A1=>
      max_calc_comparator_fourth_inp1_8, B0=>nx15492, B1=>nx15730);
   max_calc_reg_comparator_fourth_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx32319, D=>nx23463, CLK=>clk);
   ix23464 : oai21 port map ( Y=>nx23463, A0=>nx32319, A1=>nx34791, B0=>
      nx32322);
   ix23474 : oai21 port map ( Y=>nx23473, A0=>nx32326, A1=>nx34793, B0=>
      nx32328);
   max_calc_reg_comparator_fourth_inp1_8 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_8, QB=>nx32326, D=>nx23473, CLK=>clk);
   ix15731 : oai22 port map ( Y=>nx15730, A0=>nx32332, A1=>nx32345, B0=>
      max_calc_comparator_fourth_inp2_7, B1=>nx32340);
   ix23484 : oai21 port map ( Y=>nx23483, A0=>nx32336, A1=>nx34793, B0=>
      nx32338);
   max_calc_reg_comparator_fourth_inp2_7 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_7, QB=>nx32336, D=>nx23483, CLK=>clk);
   ix32339 : nand03 port map ( Y=>nx32338, A0=>label_8_output(7), A1=>
      nx35465, A2=>nx34793);
   max_calc_reg_comparator_fourth_inp1_7 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_7, QB=>nx32340, D=>nx23493, CLK=>clk);
   ix23494 : oai21 port map ( Y=>nx23493, A0=>nx32340, A1=>nx34793, B0=>
      nx32343);
   ix32344 : nand03 port map ( Y=>nx32343, A0=>label_7_output(7), A1=>
      nx35467, A2=>nx34793);
   ix32346 : aoi22 port map ( Y=>nx32345, A0=>nx32347, A1=>
      max_calc_comparator_fourth_inp1_6, B0=>nx15536, B1=>nx15714);
   max_calc_reg_comparator_fourth_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx32347, D=>nx23503, CLK=>clk);
   ix23504 : oai21 port map ( Y=>nx23503, A0=>nx32347, A1=>nx34793, B0=>
      nx32350);
   ix23514 : oai21 port map ( Y=>nx23513, A0=>nx32354, A1=>nx34795, B0=>
      nx32356);
   max_calc_reg_comparator_fourth_inp1_6 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_6, QB=>nx32354, D=>nx23513, CLK=>clk);
   ix15715 : oai22 port map ( Y=>nx15714, A0=>nx32360, A1=>nx32373, B0=>
      max_calc_comparator_fourth_inp2_5, B1=>nx32368);
   ix23524 : oai21 port map ( Y=>nx23523, A0=>nx32364, A1=>nx34795, B0=>
      nx32366);
   max_calc_reg_comparator_fourth_inp2_5 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_5, QB=>nx32364, D=>nx23523, CLK=>clk);
   ix32367 : nand03 port map ( Y=>nx32366, A0=>label_8_output(5), A1=>
      nx35467, A2=>nx34795);
   max_calc_reg_comparator_fourth_inp1_5 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_5, QB=>nx32368, D=>nx23533, CLK=>clk);
   ix23534 : oai21 port map ( Y=>nx23533, A0=>nx32368, A1=>nx34795, B0=>
      nx32371);
   ix32372 : nand03 port map ( Y=>nx32371, A0=>label_7_output(5), A1=>
      nx35467, A2=>nx34795);
   ix32374 : aoi22 port map ( Y=>nx32373, A0=>nx32375, A1=>
      max_calc_comparator_fourth_inp1_4, B0=>nx15580, B1=>nx15698);
   max_calc_reg_comparator_fourth_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx32375, D=>nx23543, CLK=>clk);
   ix23544 : oai21 port map ( Y=>nx23543, A0=>nx32375, A1=>nx34797, B0=>
      nx32378);
   ix23554 : oai21 port map ( Y=>nx23553, A0=>nx32382, A1=>nx34797, B0=>
      nx32384);
   max_calc_reg_comparator_fourth_inp1_4 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_4, QB=>nx32382, D=>nx23553, CLK=>clk);
   ix15699 : oai22 port map ( Y=>nx15698, A0=>nx32388, A1=>nx32401, B0=>
      max_calc_comparator_fourth_inp2_3, B1=>nx32396);
   ix23564 : oai21 port map ( Y=>nx23563, A0=>nx32392, A1=>nx34797, B0=>
      nx32394);
   max_calc_reg_comparator_fourth_inp2_3 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_3, QB=>nx32392, D=>nx23563, CLK=>clk);
   ix32395 : nand03 port map ( Y=>nx32394, A0=>label_8_output(3), A1=>
      nx35469, A2=>nx34797);
   max_calc_reg_comparator_fourth_inp1_3 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_3, QB=>nx32396, D=>nx23573, CLK=>clk);
   ix23574 : oai21 port map ( Y=>nx23573, A0=>nx32396, A1=>nx34797, B0=>
      nx32399);
   ix32400 : nand03 port map ( Y=>nx32399, A0=>label_7_output(3), A1=>
      nx35469, A2=>nx34799);
   ix32402 : aoi22 port map ( Y=>nx32401, A0=>nx32403, A1=>
      max_calc_comparator_fourth_inp1_2, B0=>nx15624, B1=>nx15682);
   max_calc_reg_comparator_fourth_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx32403, D=>nx23583, CLK=>clk);
   ix23584 : oai21 port map ( Y=>nx23583, A0=>nx32403, A1=>nx34799, B0=>
      nx32406);
   ix23594 : oai21 port map ( Y=>nx23593, A0=>nx32410, A1=>nx34799, B0=>
      nx32412);
   max_calc_reg_comparator_fourth_inp1_2 : dff port map ( Q=>
      max_calc_comparator_fourth_inp1_2, QB=>nx32410, D=>nx23593, CLK=>clk);
   ix15683 : oai21 port map ( Y=>nx15682, A0=>
      max_calc_comparator_fourth_inp2_1, A1=>nx32422, B0=>nx32427);
   ix23604 : oai21 port map ( Y=>nx23603, A0=>nx32418, A1=>nx34799, B0=>
      nx32420);
   max_calc_reg_comparator_fourth_inp2_1 : dff port map ( Q=>
      max_calc_comparator_fourth_inp2_1, QB=>nx32418, D=>nx23603, CLK=>clk);
   ix32421 : nand03 port map ( Y=>nx32420, A0=>label_8_output(1), A1=>
      nx35469, A2=>nx34799);
   max_calc_reg_comparator_fourth_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx32422, D=>nx23613, CLK=>clk);
   ix23614 : oai21 port map ( Y=>nx23613, A0=>nx32422, A1=>nx34801, B0=>
      nx32425);
   ix32426 : nand03 port map ( Y=>nx32425, A0=>label_7_output(1), A1=>
      nx35469, A2=>nx34801);
   ix32428 : oai21 port map ( Y=>nx32427, A0=>nx31429, A1=>
      max_calc_comparator_fourth_inp1_0, B0=>nx15646);
   ix23664 : oai21 port map ( Y=>nx23663, A0=>nx32433, A1=>nx34801, B0=>
      nx32435);
   max_calc_reg_comparator_fourth_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx32433, D=>nx23663, CLK=>clk);
   ix32436 : nand03 port map ( Y=>nx32435, A0=>label_8_output(15), A1=>
      nx35469, A2=>nx34801);
   labelsregfile_label8_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_8_output(15), QB=>OPEN, D=>nx23653, CLK=>clk, R=>rst);
   lat_label_8_input_15 : latch port map ( Q=>label_8_input_15, D=>nx15808, 
      CLK=>nx34539);
   reg_label_8_input_state_machine_15 : dffr port map ( Q=>
      label_8_input_state_machine_15, QB=>OPEN, D=>nx23643, CLK=>clk, R=>rst
   );
   ix15805 : xnor2 port map ( Y=>nx15804, A0=>nx15800, A1=>nx32446);
   ix15801 : oai22 port map ( Y=>nx15800, A0=>nx31882, A1=>nx32054, B0=>
      nx32056, B1=>nx31850);
   ix23694 : oai21 port map ( Y=>nx23693, A0=>nx32451, A1=>nx34801, B0=>
      nx32453);
   max_calc_reg_comparator_fourth_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx32451, D=>nx23693, CLK=>clk);
   labelsregfile_label7_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_7_output(15), QB=>OPEN, D=>nx23683, CLK=>clk, R=>rst);
   lat_label_7_input_15 : latch port map ( Q=>label_7_input_15, D=>nx15850, 
      CLK=>nx34539);
   reg_label_7_input_state_machine_15 : dffr port map ( Q=>
      label_7_input_state_machine_15, QB=>OPEN, D=>nx23673, CLK=>clk, R=>rst
   );
   ix15847 : xnor2 port map ( Y=>nx15846, A0=>nx15842, A1=>nx32464);
   ix15843 : oai22 port map ( Y=>nx15842, A0=>nx32071, A1=>nx32243, B0=>
      nx32245, B1=>nx31411);
   max_calc_reg_ans4_0 : dff port map ( Q=>max_calc_ans4_0, QB=>OPEN, D=>
      nx24243, CLK=>clk);
   ix17139 : xnor2 port map ( Y=>nx17138, A0=>nx32470, A1=>nx17136);
   ix32471 : aoi22 port map ( Y=>nx32470, A0=>nx32472, A1=>
      max_calc_comparator_second_inp1_14, B0=>nx15908, B1=>nx17054);
   max_calc_reg_comparator_second_inp2_14 : dff port map ( Q=>OPEN, QB=>
      nx32472, D=>nx23713, CLK=>clk);
   ix23714 : oai21 port map ( Y=>nx23713, A0=>nx32472, A1=>nx34803, B0=>
      nx32475);
   ix32476 : nand03 port map ( Y=>nx32475, A0=>nx35175, A1=>nx15896, A2=>
      nx34803);
   labelsregfile_label4_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_4_output(14), QB=>nx32660, D=>nx14953, CLK=>clk, R=>rst);
   lat_label_4_input_14 : latch port map ( Q=>label_4_input_14, D=>nx2186, 
      CLK=>nx34543);
   reg_label_4_input_state_machine_14 : dffr port map ( Q=>
      label_4_input_state_machine_14, QB=>OPEN, D=>nx14943, CLK=>clk, R=>rst
   );
   ix2183 : xor2 port map ( Y=>nx2182, A0=>nx32486, A1=>nx32658);
   ix32487 : aoi22 port map ( Y=>nx32486, A0=>label_4_output(13), A1=>
      booth_booth_integration_output_3_13, B0=>nx2140, B1=>nx12959);
   labelsregfile_label4_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_4_output(13), QB=>OPEN, D=>nx14933, CLK=>clk, R=>rst);
   lat_label_4_input_13 : latch port map ( Q=>label_4_input_13, D=>nx2154, 
      CLK=>nx34543);
   reg_label_4_input_state_machine_13 : dffr port map ( Q=>
      label_4_input_state_machine_13, QB=>OPEN, D=>nx14923, CLK=>clk, R=>rst
   );
   ix2151 : xnor2 port map ( Y=>nx2150, A0=>nx2140, A1=>nx32654);
   ix2141 : oai22 port map ( Y=>nx2140, A0=>nx32497, A1=>nx32643, B0=>
      nx32653, B1=>nx30970);
   ix32498 : aoi22 port map ( Y=>nx32497, A0=>label_4_output(11), A1=>
      booth_booth_integration_output_3_11, B0=>nx2076, B1=>nx12955);
   labelsregfile_label4_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_4_output(11), QB=>OPEN, D=>nx14893, CLK=>clk, R=>rst);
   lat_label_4_input_11 : latch port map ( Q=>label_4_input_11, D=>nx2090, 
      CLK=>nx34541);
   reg_label_4_input_state_machine_11 : dffr port map ( Q=>
      label_4_input_state_machine_11, QB=>OPEN, D=>nx14883, CLK=>clk, R=>rst
   );
   ix2087 : xnor2 port map ( Y=>nx2086, A0=>nx2076, A1=>nx32639);
   ix2077 : oai22 port map ( Y=>nx2076, A0=>nx32508, A1=>nx32628, B0=>
      nx32638, B1=>nx30972);
   ix32509 : aoi22 port map ( Y=>nx32508, A0=>label_4_output(9), A1=>
      booth_booth_integration_output_3_9, B0=>nx2012, B1=>nx12953);
   labelsregfile_label4_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_4_output(9), QB=>OPEN, D=>nx14853, CLK=>clk, R=>rst);
   lat_label_4_input_9 : latch port map ( Q=>label_4_input_9, D=>nx2026, CLK
      =>nx34541);
   reg_label_4_input_state_machine_9 : dffr port map ( Q=>
      label_4_input_state_machine_9, QB=>OPEN, D=>nx14843, CLK=>clk, R=>rst
   );
   ix2023 : xnor2 port map ( Y=>nx2022, A0=>nx2012, A1=>nx32624);
   ix2013 : oai22 port map ( Y=>nx2012, A0=>nx32519, A1=>nx32613, B0=>
      nx32623, B1=>nx30974);
   ix32520 : aoi22 port map ( Y=>nx32519, A0=>label_4_output(7), A1=>
      booth_booth_integration_output_3_7, B0=>nx1948, B1=>nx12949);
   labelsregfile_label4_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_4_output(7), QB=>OPEN, D=>nx14813, CLK=>clk, R=>rst);
   lat_label_4_input_7 : latch port map ( Q=>label_4_input_7, D=>nx1962, CLK
      =>nx34541);
   reg_label_4_input_state_machine_7 : dffr port map ( Q=>
      label_4_input_state_machine_7, QB=>OPEN, D=>nx14803, CLK=>clk, R=>rst
   );
   ix1959 : xnor2 port map ( Y=>nx1958, A0=>nx1948, A1=>nx32609);
   ix1949 : oai22 port map ( Y=>nx1948, A0=>nx32530, A1=>nx32598, B0=>
      nx32608, B1=>nx30976);
   ix32531 : aoi22 port map ( Y=>nx32530, A0=>label_4_output(5), A1=>
      booth_booth_integration_output_3_5, B0=>nx1884, B1=>nx12946);
   labelsregfile_label4_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_4_output(5), QB=>OPEN, D=>nx14773, CLK=>clk, R=>rst);
   lat_label_4_input_5 : latch port map ( Q=>label_4_input_5, D=>nx1898, CLK
      =>nx34539);
   reg_label_4_input_state_machine_5 : dffr port map ( Q=>
      label_4_input_state_machine_5, QB=>OPEN, D=>nx14763, CLK=>clk, R=>rst
   );
   ix1895 : xnor2 port map ( Y=>nx1894, A0=>nx1884, A1=>nx32594);
   ix1885 : oai22 port map ( Y=>nx1884, A0=>nx32541, A1=>nx32583, B0=>
      nx32593, B1=>nx30978);
   ix32542 : aoi22 port map ( Y=>nx32541, A0=>label_4_output(3), A1=>
      booth_booth_integration_output_3_3, B0=>nx1820, B1=>nx12943);
   labelsregfile_label4_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_4_output(3), QB=>OPEN, D=>nx14733, CLK=>clk, R=>rst);
   lat_label_4_input_3 : latch port map ( Q=>label_4_input_3, D=>nx1834, CLK
      =>nx34539);
   reg_label_4_input_state_machine_3 : dffr port map ( Q=>
      label_4_input_state_machine_3, QB=>OPEN, D=>nx14723, CLK=>clk, R=>rst
   );
   ix1831 : xnor2 port map ( Y=>nx1830, A0=>nx1820, A1=>nx32579);
   ix1821 : oai22 port map ( Y=>nx1820, A0=>nx32552, A1=>nx32568, B0=>
      nx32578, B1=>nx30980);
   ix32553 : aoi32 port map ( Y=>nx32552, A0=>label_4_output(0), A1=>nx35719, 
      A2=>nx12939, B0=>label_4_output(1), B1=>
      booth_booth_integration_output_3_1);
   labelsregfile_label4_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_4_output(1), QB=>OPEN, D=>nx14693, CLK=>clk, R=>rst);
   lat_label_4_input_1 : latch port map ( Q=>label_4_input_1, D=>nx1770, CLK
      =>nx34539);
   reg_label_4_input_state_machine_1 : dffr port map ( Q=>
      label_4_input_state_machine_1, QB=>OPEN, D=>nx14683, CLK=>clk, R=>rst
   );
   ix1767 : xor2 port map ( Y=>nx1766, A0=>nx32563, A1=>nx32565);
   ix32564 : nand02 port map ( Y=>nx32563, A0=>label_4_output(0), A1=>
      nx35719);
   ix32566 : xnor2 port map ( Y=>nx32565, A0=>
      booth_booth_integration_output_3_1, A1=>label_4_output(1));
   labelsregfile_label4_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_4_output(2), QB=>nx32578, D=>nx14713, CLK=>clk, R=>rst);
   lat_label_4_input_2 : latch port map ( Q=>label_4_input_2, D=>nx1802, CLK
      =>nx34539);
   reg_label_4_input_state_machine_2 : dffr port map ( Q=>
      label_4_input_state_machine_2, QB=>OPEN, D=>nx14703, CLK=>clk, R=>rst
   );
   ix1799 : xor2 port map ( Y=>nx1798, A0=>nx32552, A1=>nx32568);
   ix32580 : xnor2 port map ( Y=>nx32579, A0=>
      booth_booth_integration_output_3_3, A1=>label_4_output(3));
   labelsregfile_label4_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_4_output(4), QB=>nx32593, D=>nx14753, CLK=>clk, R=>rst);
   lat_label_4_input_4 : latch port map ( Q=>label_4_input_4, D=>nx1866, CLK
      =>nx34539);
   reg_label_4_input_state_machine_4 : dffr port map ( Q=>
      label_4_input_state_machine_4, QB=>OPEN, D=>nx14743, CLK=>clk, R=>rst
   );
   ix1863 : xor2 port map ( Y=>nx1862, A0=>nx32541, A1=>nx32583);
   ix32595 : xnor2 port map ( Y=>nx32594, A0=>
      booth_booth_integration_output_3_5, A1=>label_4_output(5));
   labelsregfile_label4_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_4_output(6), QB=>nx32608, D=>nx14793, CLK=>clk, R=>rst);
   lat_label_4_input_6 : latch port map ( Q=>label_4_input_6, D=>nx1930, CLK
      =>nx34541);
   reg_label_4_input_state_machine_6 : dffr port map ( Q=>
      label_4_input_state_machine_6, QB=>OPEN, D=>nx14783, CLK=>clk, R=>rst
   );
   ix1927 : xor2 port map ( Y=>nx1926, A0=>nx32530, A1=>nx32598);
   ix32610 : xnor2 port map ( Y=>nx32609, A0=>
      booth_booth_integration_output_3_7, A1=>label_4_output(7));
   labelsregfile_label4_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_4_output(8), QB=>nx32623, D=>nx14833, CLK=>clk, R=>rst);
   lat_label_4_input_8 : latch port map ( Q=>label_4_input_8, D=>nx1994, CLK
      =>nx34541);
   reg_label_4_input_state_machine_8 : dffr port map ( Q=>
      label_4_input_state_machine_8, QB=>OPEN, D=>nx14823, CLK=>clk, R=>rst
   );
   ix1991 : xor2 port map ( Y=>nx1990, A0=>nx32519, A1=>nx32613);
   ix32625 : xnor2 port map ( Y=>nx32624, A0=>
      booth_booth_integration_output_3_9, A1=>label_4_output(9));
   labelsregfile_label4_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_4_output(10), QB=>nx32638, D=>nx14873, CLK=>clk, R=>rst);
   lat_label_4_input_10 : latch port map ( Q=>label_4_input_10, D=>nx2058, 
      CLK=>nx34541);
   reg_label_4_input_state_machine_10 : dffr port map ( Q=>
      label_4_input_state_machine_10, QB=>OPEN, D=>nx14863, CLK=>clk, R=>rst
   );
   ix2055 : xor2 port map ( Y=>nx2054, A0=>nx32508, A1=>nx32628);
   ix32640 : xnor2 port map ( Y=>nx32639, A0=>
      booth_booth_integration_output_3_11, A1=>label_4_output(11));
   labelsregfile_label4_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_4_output(12), QB=>nx32653, D=>nx14913, CLK=>clk, R=>rst);
   lat_label_4_input_12 : latch port map ( Q=>label_4_input_12, D=>nx2122, 
      CLK=>nx34541);
   reg_label_4_input_state_machine_12 : dffr port map ( Q=>
      label_4_input_state_machine_12, QB=>OPEN, D=>nx14903, CLK=>clk, R=>rst
   );
   ix2119 : xor2 port map ( Y=>nx2118, A0=>nx32497, A1=>nx32643);
   ix32655 : xnor2 port map ( Y=>nx32654, A0=>
      booth_booth_integration_output_3_13, A1=>label_4_output(13));
   max_calc_reg_ans4_14 : dff port map ( Q=>max_calc_ans4_14, QB=>nx32665, D
      =>nx23703, CLK=>clk);
   ix21674 : oai21 port map ( Y=>nx21673, A0=>nx32669, A1=>nx34803, B0=>
      nx32671);
   max_calc_reg_comparator_second_inp1_14 : dff port map ( Q=>
      max_calc_comparator_second_inp1_14, QB=>nx32669, D=>nx21673, CLK=>clk
   );
   ix32672 : nand03 port map ( Y=>nx32671, A0=>nx35175, A1=>nx12712, A2=>
      nx34803);
   labelsregfile_label3_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_3_output(14), QB=>nx32856, D=>nx15803, CLK=>clk, R=>rst);
   lat_label_3_input_14 : latch port map ( Q=>label_3_input_14, D=>nx3524, 
      CLK=>nx34547);
   reg_label_3_input_state_machine_14 : dffr port map ( Q=>
      label_3_input_state_machine_14, QB=>OPEN, D=>nx15793, CLK=>clk, R=>rst
   );
   ix3521 : xor2 port map ( Y=>nx3520, A0=>nx32682, A1=>nx32854);
   ix32683 : aoi22 port map ( Y=>nx32682, A0=>label_3_output(13), A1=>
      booth_booth_integration_output_2_13, B0=>nx3478, B1=>nx13011);
   labelsregfile_label3_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_3_output(13), QB=>OPEN, D=>nx15783, CLK=>clk, R=>rst);
   lat_label_3_input_13 : latch port map ( Q=>label_3_input_13, D=>nx3492, 
      CLK=>nx34547);
   reg_label_3_input_state_machine_13 : dffr port map ( Q=>
      label_3_input_state_machine_13, QB=>OPEN, D=>nx15773, CLK=>clk, R=>rst
   );
   ix3489 : xnor2 port map ( Y=>nx3488, A0=>nx3478, A1=>nx32850);
   ix3479 : oai22 port map ( Y=>nx3478, A0=>nx32693, A1=>nx32839, B0=>
      nx32849, B1=>nx29041);
   ix32694 : aoi22 port map ( Y=>nx32693, A0=>label_3_output(11), A1=>
      booth_booth_integration_output_2_11, B0=>nx3414, B1=>nx13007);
   labelsregfile_label3_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_3_output(11), QB=>OPEN, D=>nx15743, CLK=>clk, R=>rst);
   lat_label_3_input_11 : latch port map ( Q=>label_3_input_11, D=>nx3428, 
      CLK=>nx34545);
   reg_label_3_input_state_machine_11 : dffr port map ( Q=>
      label_3_input_state_machine_11, QB=>OPEN, D=>nx15733, CLK=>clk, R=>rst
   );
   ix3425 : xnor2 port map ( Y=>nx3424, A0=>nx3414, A1=>nx32835);
   ix3415 : oai22 port map ( Y=>nx3414, A0=>nx32704, A1=>nx32824, B0=>
      nx32834, B1=>nx29043);
   ix32705 : aoi22 port map ( Y=>nx32704, A0=>label_3_output(9), A1=>
      booth_booth_integration_output_2_9, B0=>nx3350, B1=>nx13003);
   labelsregfile_label3_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_3_output(9), QB=>OPEN, D=>nx15703, CLK=>clk, R=>rst);
   lat_label_3_input_9 : latch port map ( Q=>label_3_input_9, D=>nx3364, CLK
      =>nx34545);
   reg_label_3_input_state_machine_9 : dffr port map ( Q=>
      label_3_input_state_machine_9, QB=>OPEN, D=>nx15693, CLK=>clk, R=>rst
   );
   ix3361 : xnor2 port map ( Y=>nx3360, A0=>nx3350, A1=>nx32820);
   ix3351 : oai22 port map ( Y=>nx3350, A0=>nx32715, A1=>nx32809, B0=>
      nx32819, B1=>nx29045);
   ix32716 : aoi22 port map ( Y=>nx32715, A0=>label_3_output(7), A1=>
      booth_booth_integration_output_2_7, B0=>nx3286, B1=>nx13001);
   labelsregfile_label3_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_3_output(7), QB=>OPEN, D=>nx15663, CLK=>clk, R=>rst);
   lat_label_3_input_7 : latch port map ( Q=>label_3_input_7, D=>nx3300, CLK
      =>nx34545);
   reg_label_3_input_state_machine_7 : dffr port map ( Q=>
      label_3_input_state_machine_7, QB=>OPEN, D=>nx15653, CLK=>clk, R=>rst
   );
   ix3297 : xnor2 port map ( Y=>nx3296, A0=>nx3286, A1=>nx32805);
   ix3287 : oai22 port map ( Y=>nx3286, A0=>nx32726, A1=>nx32794, B0=>
      nx32804, B1=>nx29047);
   ix32727 : aoi22 port map ( Y=>nx32726, A0=>label_3_output(5), A1=>
      booth_booth_integration_output_2_5, B0=>nx3222, B1=>nx12997);
   labelsregfile_label3_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_3_output(5), QB=>OPEN, D=>nx15623, CLK=>clk, R=>rst);
   lat_label_3_input_5 : latch port map ( Q=>label_3_input_5, D=>nx3236, CLK
      =>nx34543);
   reg_label_3_input_state_machine_5 : dffr port map ( Q=>
      label_3_input_state_machine_5, QB=>OPEN, D=>nx15613, CLK=>clk, R=>rst
   );
   ix3233 : xnor2 port map ( Y=>nx3232, A0=>nx3222, A1=>nx32790);
   ix3223 : oai22 port map ( Y=>nx3222, A0=>nx32737, A1=>nx32779, B0=>
      nx32789, B1=>nx29049);
   ix32738 : aoi22 port map ( Y=>nx32737, A0=>label_3_output(3), A1=>
      booth_booth_integration_output_2_3, B0=>nx3158, B1=>nx12994);
   labelsregfile_label3_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_3_output(3), QB=>OPEN, D=>nx15583, CLK=>clk, R=>rst);
   lat_label_3_input_3 : latch port map ( Q=>label_3_input_3, D=>nx3172, CLK
      =>nx34543);
   reg_label_3_input_state_machine_3 : dffr port map ( Q=>
      label_3_input_state_machine_3, QB=>OPEN, D=>nx15573, CLK=>clk, R=>rst
   );
   ix3169 : xnor2 port map ( Y=>nx3168, A0=>nx3158, A1=>nx32775);
   ix3159 : oai22 port map ( Y=>nx3158, A0=>nx32748, A1=>nx32764, B0=>
      nx32774, B1=>nx29051);
   ix32749 : aoi32 port map ( Y=>nx32748, A0=>label_3_output(0), A1=>nx35723, 
      A2=>nx12991, B0=>label_3_output(1), B1=>
      booth_booth_integration_output_2_1);
   labelsregfile_label3_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_3_output(1), QB=>OPEN, D=>nx15543, CLK=>clk, R=>rst);
   lat_label_3_input_1 : latch port map ( Q=>label_3_input_1, D=>nx3108, CLK
      =>nx34543);
   reg_label_3_input_state_machine_1 : dffr port map ( Q=>
      label_3_input_state_machine_1, QB=>OPEN, D=>nx15533, CLK=>clk, R=>rst
   );
   ix3105 : xor2 port map ( Y=>nx3104, A0=>nx32759, A1=>nx32761);
   ix32760 : nand02 port map ( Y=>nx32759, A0=>label_3_output(0), A1=>
      nx35723);
   ix32762 : xnor2 port map ( Y=>nx32761, A0=>
      booth_booth_integration_output_2_1, A1=>label_3_output(1));
   labelsregfile_label3_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_3_output(2), QB=>nx32774, D=>nx15563, CLK=>clk, R=>rst);
   lat_label_3_input_2 : latch port map ( Q=>label_3_input_2, D=>nx3140, CLK
      =>nx34543);
   reg_label_3_input_state_machine_2 : dffr port map ( Q=>
      label_3_input_state_machine_2, QB=>OPEN, D=>nx15553, CLK=>clk, R=>rst
   );
   ix3137 : xor2 port map ( Y=>nx3136, A0=>nx32748, A1=>nx32764);
   ix32776 : xnor2 port map ( Y=>nx32775, A0=>
      booth_booth_integration_output_2_3, A1=>label_3_output(3));
   labelsregfile_label3_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_3_output(4), QB=>nx32789, D=>nx15603, CLK=>clk, R=>rst);
   lat_label_3_input_4 : latch port map ( Q=>label_3_input_4, D=>nx3204, CLK
      =>nx34543);
   reg_label_3_input_state_machine_4 : dffr port map ( Q=>
      label_3_input_state_machine_4, QB=>OPEN, D=>nx15593, CLK=>clk, R=>rst
   );
   ix3201 : xor2 port map ( Y=>nx3200, A0=>nx32737, A1=>nx32779);
   ix32791 : xnor2 port map ( Y=>nx32790, A0=>
      booth_booth_integration_output_2_5, A1=>label_3_output(5));
   labelsregfile_label3_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_3_output(6), QB=>nx32804, D=>nx15643, CLK=>clk, R=>rst);
   lat_label_3_input_6 : latch port map ( Q=>label_3_input_6, D=>nx3268, CLK
      =>nx34545);
   reg_label_3_input_state_machine_6 : dffr port map ( Q=>
      label_3_input_state_machine_6, QB=>OPEN, D=>nx15633, CLK=>clk, R=>rst
   );
   ix3265 : xor2 port map ( Y=>nx3264, A0=>nx32726, A1=>nx32794);
   ix32806 : xnor2 port map ( Y=>nx32805, A0=>
      booth_booth_integration_output_2_7, A1=>label_3_output(7));
   labelsregfile_label3_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_3_output(8), QB=>nx32819, D=>nx15683, CLK=>clk, R=>rst);
   lat_label_3_input_8 : latch port map ( Q=>label_3_input_8, D=>nx3332, CLK
      =>nx34545);
   reg_label_3_input_state_machine_8 : dffr port map ( Q=>
      label_3_input_state_machine_8, QB=>OPEN, D=>nx15673, CLK=>clk, R=>rst
   );
   ix3329 : xor2 port map ( Y=>nx3328, A0=>nx32715, A1=>nx32809);
   ix32821 : xnor2 port map ( Y=>nx32820, A0=>
      booth_booth_integration_output_2_9, A1=>label_3_output(9));
   labelsregfile_label3_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_3_output(10), QB=>nx32834, D=>nx15723, CLK=>clk, R=>rst);
   lat_label_3_input_10 : latch port map ( Q=>label_3_input_10, D=>nx3396, 
      CLK=>nx34545);
   reg_label_3_input_state_machine_10 : dffr port map ( Q=>
      label_3_input_state_machine_10, QB=>OPEN, D=>nx15713, CLK=>clk, R=>rst
   );
   ix3393 : xor2 port map ( Y=>nx3392, A0=>nx32704, A1=>nx32824);
   ix32836 : xnor2 port map ( Y=>nx32835, A0=>
      booth_booth_integration_output_2_11, A1=>label_3_output(11));
   labelsregfile_label3_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_3_output(12), QB=>nx32849, D=>nx15763, CLK=>clk, R=>rst);
   lat_label_3_input_12 : latch port map ( Q=>label_3_input_12, D=>nx3460, 
      CLK=>nx34545);
   reg_label_3_input_state_machine_12 : dffr port map ( Q=>
      label_3_input_state_machine_12, QB=>OPEN, D=>nx15753, CLK=>clk, R=>rst
   );
   ix3457 : xor2 port map ( Y=>nx3456, A0=>nx32693, A1=>nx32839);
   ix32851 : xnor2 port map ( Y=>nx32850, A0=>
      booth_booth_integration_output_2_13, A1=>label_3_output(13));
   max_calc_reg_ans3_14 : dff port map ( Q=>max_calc_ans3_14, QB=>nx32861, D
      =>nx21663, CLK=>clk);
   ix17055 : oai22 port map ( Y=>nx17054, A0=>nx32865, A1=>nx32892, B0=>
      max_calc_comparator_second_inp2_13, B1=>nx32880);
   ix23734 : oai21 port map ( Y=>nx23733, A0=>nx32869, A1=>nx34803, B0=>
      nx32871);
   max_calc_reg_comparator_second_inp2_13 : dff port map ( Q=>
      max_calc_comparator_second_inp2_13, QB=>nx32869, D=>nx23733, CLK=>clk
   );
   ix32872 : nand03 port map ( Y=>nx32871, A0=>nx35175, A1=>nx15934, A2=>
      nx34803);
   max_calc_reg_ans4_13 : dff port map ( Q=>max_calc_ans4_13, QB=>OPEN, D=>
      nx23723, CLK=>clk);
   max_calc_reg_comparator_second_inp1_13 : dff port map ( Q=>
      max_calc_comparator_second_inp1_13, QB=>nx32880, D=>nx23753, CLK=>clk
   );
   ix23754 : oai21 port map ( Y=>nx23753, A0=>nx32880, A1=>nx34803, B0=>
      nx32883);
   ix32884 : nand03 port map ( Y=>nx32883, A0=>nx35175, A1=>nx15970, A2=>
      nx34805);
   max_calc_reg_ans3_13 : dff port map ( Q=>max_calc_ans3_13, QB=>OPEN, D=>
      nx23743, CLK=>clk);
   ix32893 : aoi22 port map ( Y=>nx32892, A0=>nx32894, A1=>
      max_calc_comparator_second_inp1_12, B0=>nx16056, B1=>nx17038);
   max_calc_reg_comparator_second_inp2_12 : dff port map ( Q=>OPEN, QB=>
      nx32894, D=>nx23773, CLK=>clk);
   ix23774 : oai21 port map ( Y=>nx23773, A0=>nx32894, A1=>nx34805, B0=>
      nx32897);
   ix32898 : nand03 port map ( Y=>nx32897, A0=>nx35175, A1=>nx16008, A2=>
      nx34805);
   max_calc_reg_ans4_12 : dff port map ( Q=>max_calc_ans4_12, QB=>nx32904, D
      =>nx23763, CLK=>clk);
   ix23794 : oai21 port map ( Y=>nx23793, A0=>nx32908, A1=>nx34805, B0=>
      nx32910);
   max_calc_reg_comparator_second_inp1_12 : dff port map ( Q=>
      max_calc_comparator_second_inp1_12, QB=>nx32908, D=>nx23793, CLK=>clk
   );
   ix32911 : nand03 port map ( Y=>nx32910, A0=>nx35175, A1=>nx16044, A2=>
      nx34805);
   max_calc_reg_ans3_12 : dff port map ( Q=>max_calc_ans3_12, QB=>nx32917, D
      =>nx23783, CLK=>clk);
   ix17039 : oai22 port map ( Y=>nx17038, A0=>nx32921, A1=>nx32948, B0=>
      max_calc_comparator_second_inp2_11, B1=>nx32936);
   ix23814 : oai21 port map ( Y=>nx23813, A0=>nx32925, A1=>nx34805, B0=>
      nx32927);
   max_calc_reg_comparator_second_inp2_11 : dff port map ( Q=>
      max_calc_comparator_second_inp2_11, QB=>nx32925, D=>nx23813, CLK=>clk
   );
   ix32928 : nand03 port map ( Y=>nx32927, A0=>nx35177, A1=>nx16082, A2=>
      nx34805);
   max_calc_reg_ans4_11 : dff port map ( Q=>max_calc_ans4_11, QB=>OPEN, D=>
      nx23803, CLK=>clk);
   max_calc_reg_comparator_second_inp1_11 : dff port map ( Q=>
      max_calc_comparator_second_inp1_11, QB=>nx32936, D=>nx23833, CLK=>clk
   );
   ix23834 : oai21 port map ( Y=>nx23833, A0=>nx32936, A1=>nx34807, B0=>
      nx32939);
   ix32940 : nand03 port map ( Y=>nx32939, A0=>nx35177, A1=>nx16118, A2=>
      nx34807);
   max_calc_reg_ans3_11 : dff port map ( Q=>max_calc_ans3_11, QB=>OPEN, D=>
      nx23823, CLK=>clk);
   ix32949 : aoi22 port map ( Y=>nx32948, A0=>nx32950, A1=>
      max_calc_comparator_second_inp1_10, B0=>nx16204, B1=>nx17022);
   max_calc_reg_comparator_second_inp2_10 : dff port map ( Q=>OPEN, QB=>
      nx32950, D=>nx23853, CLK=>clk);
   ix23854 : oai21 port map ( Y=>nx23853, A0=>nx32950, A1=>nx34807, B0=>
      nx32953);
   ix32954 : nand03 port map ( Y=>nx32953, A0=>nx35177, A1=>nx16156, A2=>
      nx34807);
   max_calc_reg_ans4_10 : dff port map ( Q=>max_calc_ans4_10, QB=>nx32960, D
      =>nx23843, CLK=>clk);
   ix23874 : oai21 port map ( Y=>nx23873, A0=>nx32964, A1=>nx34807, B0=>
      nx32966);
   max_calc_reg_comparator_second_inp1_10 : dff port map ( Q=>
      max_calc_comparator_second_inp1_10, QB=>nx32964, D=>nx23873, CLK=>clk
   );
   ix32967 : nand03 port map ( Y=>nx32966, A0=>nx35177, A1=>nx16192, A2=>
      nx34807);
   max_calc_reg_ans3_10 : dff port map ( Q=>max_calc_ans3_10, QB=>nx32973, D
      =>nx23863, CLK=>clk);
   ix17023 : oai22 port map ( Y=>nx17022, A0=>nx32977, A1=>nx33004, B0=>
      max_calc_comparator_second_inp2_9, B1=>nx32992);
   ix23894 : oai21 port map ( Y=>nx23893, A0=>nx32981, A1=>nx34807, B0=>
      nx32983);
   max_calc_reg_comparator_second_inp2_9 : dff port map ( Q=>
      max_calc_comparator_second_inp2_9, QB=>nx32981, D=>nx23893, CLK=>clk);
   ix32984 : nand03 port map ( Y=>nx32983, A0=>nx35177, A1=>nx16230, A2=>
      nx34809);
   max_calc_reg_ans4_9 : dff port map ( Q=>max_calc_ans4_9, QB=>OPEN, D=>
      nx23883, CLK=>clk);
   max_calc_reg_comparator_second_inp1_9 : dff port map ( Q=>
      max_calc_comparator_second_inp1_9, QB=>nx32992, D=>nx23913, CLK=>clk);
   ix23914 : oai21 port map ( Y=>nx23913, A0=>nx32992, A1=>nx34809, B0=>
      nx32995);
   ix32996 : nand03 port map ( Y=>nx32995, A0=>nx35177, A1=>nx16266, A2=>
      nx34809);
   max_calc_reg_ans3_9 : dff port map ( Q=>max_calc_ans3_9, QB=>OPEN, D=>
      nx23903, CLK=>clk);
   ix33005 : aoi22 port map ( Y=>nx33004, A0=>nx33006, A1=>
      max_calc_comparator_second_inp1_8, B0=>nx16352, B1=>nx17006);
   max_calc_reg_comparator_second_inp2_8 : dff port map ( Q=>OPEN, QB=>
      nx33006, D=>nx23933, CLK=>clk);
   ix23934 : oai21 port map ( Y=>nx23933, A0=>nx33006, A1=>nx34809, B0=>
      nx33009);
   ix33010 : nand03 port map ( Y=>nx33009, A0=>nx35177, A1=>nx16304, A2=>
      nx34809);
   max_calc_reg_ans4_8 : dff port map ( Q=>max_calc_ans4_8, QB=>nx33016, D=>
      nx23923, CLK=>clk);
   ix23954 : oai21 port map ( Y=>nx23953, A0=>nx33020, A1=>nx34809, B0=>
      nx33022);
   max_calc_reg_comparator_second_inp1_8 : dff port map ( Q=>
      max_calc_comparator_second_inp1_8, QB=>nx33020, D=>nx23953, CLK=>clk);
   ix33023 : nand03 port map ( Y=>nx33022, A0=>nx35179, A1=>nx16340, A2=>
      nx34809);
   max_calc_reg_ans3_8 : dff port map ( Q=>max_calc_ans3_8, QB=>nx33029, D=>
      nx23943, CLK=>clk);
   ix17007 : oai22 port map ( Y=>nx17006, A0=>nx33033, A1=>nx33060, B0=>
      max_calc_comparator_second_inp2_7, B1=>nx33048);
   ix23974 : oai21 port map ( Y=>nx23973, A0=>nx33037, A1=>nx34811, B0=>
      nx33039);
   max_calc_reg_comparator_second_inp2_7 : dff port map ( Q=>
      max_calc_comparator_second_inp2_7, QB=>nx33037, D=>nx23973, CLK=>clk);
   ix33040 : nand03 port map ( Y=>nx33039, A0=>nx35179, A1=>nx16378, A2=>
      nx34811);
   max_calc_reg_ans4_7 : dff port map ( Q=>max_calc_ans4_7, QB=>OPEN, D=>
      nx23963, CLK=>clk);
   max_calc_reg_comparator_second_inp1_7 : dff port map ( Q=>
      max_calc_comparator_second_inp1_7, QB=>nx33048, D=>nx23993, CLK=>clk);
   ix23994 : oai21 port map ( Y=>nx23993, A0=>nx33048, A1=>nx34811, B0=>
      nx33051);
   ix33052 : nand03 port map ( Y=>nx33051, A0=>nx35179, A1=>nx16414, A2=>
      nx34811);
   max_calc_reg_ans3_7 : dff port map ( Q=>max_calc_ans3_7, QB=>OPEN, D=>
      nx23983, CLK=>clk);
   ix33061 : aoi22 port map ( Y=>nx33060, A0=>nx33062, A1=>
      max_calc_comparator_second_inp1_6, B0=>nx16500, B1=>nx16990);
   max_calc_reg_comparator_second_inp2_6 : dff port map ( Q=>OPEN, QB=>
      nx33062, D=>nx24013, CLK=>clk);
   ix24014 : oai21 port map ( Y=>nx24013, A0=>nx33062, A1=>nx34811, B0=>
      nx33065);
   ix33066 : nand03 port map ( Y=>nx33065, A0=>nx35179, A1=>nx16452, A2=>
      nx34811);
   max_calc_reg_ans4_6 : dff port map ( Q=>max_calc_ans4_6, QB=>nx33072, D=>
      nx24003, CLK=>clk);
   ix24034 : oai21 port map ( Y=>nx24033, A0=>nx33076, A1=>nx34811, B0=>
      nx33078);
   max_calc_reg_comparator_second_inp1_6 : dff port map ( Q=>
      max_calc_comparator_second_inp1_6, QB=>nx33076, D=>nx24033, CLK=>clk);
   ix33079 : nand03 port map ( Y=>nx33078, A0=>nx35179, A1=>nx16488, A2=>
      nx34813);
   max_calc_reg_ans3_6 : dff port map ( Q=>max_calc_ans3_6, QB=>nx33085, D=>
      nx24023, CLK=>clk);
   ix16991 : oai22 port map ( Y=>nx16990, A0=>nx33089, A1=>nx33116, B0=>
      max_calc_comparator_second_inp2_5, B1=>nx33104);
   ix24054 : oai21 port map ( Y=>nx24053, A0=>nx33093, A1=>nx34813, B0=>
      nx33095);
   max_calc_reg_comparator_second_inp2_5 : dff port map ( Q=>
      max_calc_comparator_second_inp2_5, QB=>nx33093, D=>nx24053, CLK=>clk);
   ix33096 : nand03 port map ( Y=>nx33095, A0=>nx35179, A1=>nx16526, A2=>
      nx34813);
   max_calc_reg_ans4_5 : dff port map ( Q=>max_calc_ans4_5, QB=>OPEN, D=>
      nx24043, CLK=>clk);
   max_calc_reg_comparator_second_inp1_5 : dff port map ( Q=>
      max_calc_comparator_second_inp1_5, QB=>nx33104, D=>nx24073, CLK=>clk);
   ix24074 : oai21 port map ( Y=>nx24073, A0=>nx33104, A1=>nx34813, B0=>
      nx33107);
   ix33108 : nand03 port map ( Y=>nx33107, A0=>nx35179, A1=>nx16562, A2=>
      nx34813);
   max_calc_reg_ans3_5 : dff port map ( Q=>max_calc_ans3_5, QB=>OPEN, D=>
      nx24063, CLK=>clk);
   ix33117 : aoi22 port map ( Y=>nx33116, A0=>nx33118, A1=>
      max_calc_comparator_second_inp1_4, B0=>nx16648, B1=>nx16974);
   max_calc_reg_comparator_second_inp2_4 : dff port map ( Q=>OPEN, QB=>
      nx33118, D=>nx24093, CLK=>clk);
   ix24094 : oai21 port map ( Y=>nx24093, A0=>nx33118, A1=>nx34813, B0=>
      nx33121);
   ix33122 : nand03 port map ( Y=>nx33121, A0=>nx35181, A1=>nx16600, A2=>
      nx34813);
   max_calc_reg_ans4_4 : dff port map ( Q=>max_calc_ans4_4, QB=>nx33128, D=>
      nx24083, CLK=>clk);
   ix24114 : oai21 port map ( Y=>nx24113, A0=>nx33132, A1=>nx34815, B0=>
      nx33134);
   max_calc_reg_comparator_second_inp1_4 : dff port map ( Q=>
      max_calc_comparator_second_inp1_4, QB=>nx33132, D=>nx24113, CLK=>clk);
   ix33135 : nand03 port map ( Y=>nx33134, A0=>nx35181, A1=>nx16636, A2=>
      nx34815);
   max_calc_reg_ans3_4 : dff port map ( Q=>max_calc_ans3_4, QB=>nx33141, D=>
      nx24103, CLK=>clk);
   ix16975 : oai22 port map ( Y=>nx16974, A0=>nx33145, A1=>nx33172, B0=>
      max_calc_comparator_second_inp2_3, B1=>nx33160);
   ix24134 : oai21 port map ( Y=>nx24133, A0=>nx33149, A1=>nx34815, B0=>
      nx33151);
   max_calc_reg_comparator_second_inp2_3 : dff port map ( Q=>
      max_calc_comparator_second_inp2_3, QB=>nx33149, D=>nx24133, CLK=>clk);
   ix33152 : nand03 port map ( Y=>nx33151, A0=>nx35181, A1=>nx16674, A2=>
      nx34815);
   max_calc_reg_ans4_3 : dff port map ( Q=>max_calc_ans4_3, QB=>OPEN, D=>
      nx24123, CLK=>clk);
   max_calc_reg_comparator_second_inp1_3 : dff port map ( Q=>
      max_calc_comparator_second_inp1_3, QB=>nx33160, D=>nx24153, CLK=>clk);
   ix24154 : oai21 port map ( Y=>nx24153, A0=>nx33160, A1=>nx34815, B0=>
      nx33163);
   ix33164 : nand03 port map ( Y=>nx33163, A0=>nx35181, A1=>nx16710, A2=>
      nx34815);
   max_calc_reg_ans3_3 : dff port map ( Q=>max_calc_ans3_3, QB=>OPEN, D=>
      nx24143, CLK=>clk);
   ix33173 : aoi22 port map ( Y=>nx33172, A0=>nx33174, A1=>
      max_calc_comparator_second_inp1_2, B0=>nx16796, B1=>nx16958);
   max_calc_reg_comparator_second_inp2_2 : dff port map ( Q=>OPEN, QB=>
      nx33174, D=>nx24173, CLK=>clk);
   ix24174 : oai21 port map ( Y=>nx24173, A0=>nx33174, A1=>nx34815, B0=>
      nx33177);
   ix33178 : nand03 port map ( Y=>nx33177, A0=>nx35181, A1=>nx16748, A2=>
      nx34817);
   max_calc_reg_ans4_2 : dff port map ( Q=>max_calc_ans4_2, QB=>nx33184, D=>
      nx24163, CLK=>clk);
   ix24194 : oai21 port map ( Y=>nx24193, A0=>nx33188, A1=>nx34817, B0=>
      nx33190);
   max_calc_reg_comparator_second_inp1_2 : dff port map ( Q=>
      max_calc_comparator_second_inp1_2, QB=>nx33188, D=>nx24193, CLK=>clk);
   ix33191 : nand03 port map ( Y=>nx33190, A0=>nx35181, A1=>nx16784, A2=>
      nx34817);
   max_calc_reg_ans3_2 : dff port map ( Q=>max_calc_ans3_2, QB=>nx33197, D=>
      nx24183, CLK=>clk);
   ix16959 : oai21 port map ( Y=>nx16958, A0=>
      max_calc_comparator_second_inp2_1, A1=>nx33214, B0=>nx33226);
   ix24214 : oai21 port map ( Y=>nx24213, A0=>nx33203, A1=>nx34817, B0=>
      nx33205);
   max_calc_reg_comparator_second_inp2_1 : dff port map ( Q=>
      max_calc_comparator_second_inp2_1, QB=>nx33203, D=>nx24213, CLK=>clk);
   ix33206 : nand03 port map ( Y=>nx33205, A0=>nx35181, A1=>nx16822, A2=>
      nx34817);
   max_calc_reg_ans4_1 : dff port map ( Q=>max_calc_ans4_1, QB=>OPEN, D=>
      nx24203, CLK=>clk);
   max_calc_reg_comparator_second_inp1_1 : dff port map ( Q=>OPEN, QB=>
      nx33214, D=>nx24233, CLK=>clk);
   ix24234 : oai21 port map ( Y=>nx24233, A0=>nx33214, A1=>nx34817, B0=>
      nx33217);
   ix33218 : nand03 port map ( Y=>nx33217, A0=>nx35959, A1=>nx16858, A2=>
      nx34817);
   max_calc_reg_ans3_1 : dff port map ( Q=>max_calc_ans3_1, QB=>OPEN, D=>
      nx24223, CLK=>clk);
   ix33227 : oai21 port map ( Y=>nx33226, A0=>nx30546, A1=>
      max_calc_comparator_second_inp1_0, B0=>nx16870);
   ix24294 : oai21 port map ( Y=>nx24293, A0=>nx33232, A1=>nx34819, B0=>
      nx33234);
   max_calc_reg_comparator_second_inp2_15 : dff port map ( Q=>OPEN, QB=>
      nx33232, D=>nx24293, CLK=>clk);
   ix33235 : nand03 port map ( Y=>nx33234, A0=>nx35959, A1=>nx17088, A2=>
      nx34819);
   labelsregfile_label4_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_4_output(15), QB=>OPEN, D=>nx14963, CLK=>clk, R=>rst);
   lat_label_4_input_15 : latch port map ( Q=>label_4_input_15, D=>nx2212, 
      CLK=>nx34547);
   reg_label_4_input_state_machine_15 : dffr port map ( Q=>
      label_4_input_state_machine_15, QB=>OPEN, D=>nx14123, CLK=>clk, R=>rst
   );
   ix2209 : xnor2 port map ( Y=>nx2208, A0=>nx2204, A1=>nx33246);
   ix2205 : oai22 port map ( Y=>nx2204, A0=>nx32486, A1=>nx32658, B0=>
      nx32660, B1=>nx30968);
   max_calc_reg_ans4_15 : dff port map ( Q=>max_calc_ans4_15, QB=>OPEN, D=>
      nx24283, CLK=>clk);
   ix24314 : oai21 port map ( Y=>nx24313, A0=>nx33257, A1=>nx34819, B0=>
      nx33259);
   max_calc_reg_comparator_second_inp1_15 : dff port map ( Q=>OPEN, QB=>
      nx33257, D=>nx24313, CLK=>clk);
   ix33260 : nand03 port map ( Y=>nx33259, A0=>nx35959, A1=>nx17124, A2=>
      nx34819);
   labelsregfile_label3_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_3_output(15), QB=>OPEN, D=>nx15813, CLK=>clk, R=>rst);
   lat_label_3_input_15 : latch port map ( Q=>label_3_input_15, D=>nx3550, 
      CLK=>nx34547);
   reg_label_3_input_state_machine_15 : dffr port map ( Q=>
      label_3_input_state_machine_15, QB=>OPEN, D=>nx14973, CLK=>clk, R=>rst
   );
   ix3547 : xnor2 port map ( Y=>nx3546, A0=>nx3542, A1=>nx33271);
   ix3543 : oai22 port map ( Y=>nx3542, A0=>nx32682, A1=>nx32854, B0=>
      nx32856, B1=>nx29039);
   max_calc_reg_ans3_15 : dff port map ( Q=>max_calc_ans3_15, QB=>OPEN, D=>
      nx24303, CLK=>clk);
   max_calc_reg_ans7_0 : dff port map ( Q=>max_calc_ans7_0, QB=>OPEN, D=>
      nx25463, CLK=>clk);
   max_calc_reg_ans8_0 : dff port map ( Q=>max_calc_ans8_0, QB=>OPEN, D=>
      nx25453, CLK=>clk);
   ix19143 : xnor2 port map ( Y=>nx13373, A0=>nx33290, A1=>nx19140);
   ix33291 : aoi22 port map ( Y=>nx33290, A0=>nx33292, A1=>
      max_calc_comparator_first_inp1_14, B0=>nx17256, B1=>nx19010);
   labelsregfile_label2_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_2_output(14), QB=>nx33479, D=>nx16653, CLK=>clk, R=>rst);
   lat_label_2_input_14 : latch port map ( Q=>label_2_input_14, D=>nx4862, 
      CLK=>nx34551);
   reg_label_2_input_state_machine_14 : dffr port map ( Q=>
      label_2_input_state_machine_14, QB=>OPEN, D=>nx16643, CLK=>clk, R=>rst
   );
   ix4859 : xor2 port map ( Y=>nx4858, A0=>nx33305, A1=>nx33477);
   ix33306 : aoi22 port map ( Y=>nx33305, A0=>label_2_output(13), A1=>
      booth_booth_integration_output_1_13, B0=>nx4816, B1=>nx13063);
   labelsregfile_label2_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_2_output(13), QB=>OPEN, D=>nx16633, CLK=>clk, R=>rst);
   lat_label_2_input_13 : latch port map ( Q=>label_2_input_13, D=>nx4830, 
      CLK=>nx34551);
   reg_label_2_input_state_machine_13 : dffr port map ( Q=>
      label_2_input_state_machine_13, QB=>OPEN, D=>nx16623, CLK=>clk, R=>rst
   );
   ix4827 : xnor2 port map ( Y=>nx4826, A0=>nx4816, A1=>nx33473);
   ix4817 : oai22 port map ( Y=>nx4816, A0=>nx33316, A1=>nx33462, B0=>
      nx33472, B1=>nx28598);
   ix33317 : aoi22 port map ( Y=>nx33316, A0=>label_2_output(11), A1=>
      booth_booth_integration_output_1_11, B0=>nx4752, B1=>nx13059);
   labelsregfile_label2_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_2_output(11), QB=>OPEN, D=>nx16593, CLK=>clk, R=>rst);
   lat_label_2_input_11 : latch port map ( Q=>label_2_input_11, D=>nx4766, 
      CLK=>nx34551);
   reg_label_2_input_state_machine_11 : dffr port map ( Q=>
      label_2_input_state_machine_11, QB=>OPEN, D=>nx16583, CLK=>clk, R=>rst
   );
   ix4763 : xnor2 port map ( Y=>nx4762, A0=>nx4752, A1=>nx33458);
   ix4753 : oai22 port map ( Y=>nx4752, A0=>nx33327, A1=>nx33447, B0=>
      nx33457, B1=>nx28600);
   ix33328 : aoi22 port map ( Y=>nx33327, A0=>label_2_output(9), A1=>
      booth_booth_integration_output_1_9, B0=>nx4688, B1=>nx13055);
   labelsregfile_label2_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_2_output(9), QB=>OPEN, D=>nx16553, CLK=>clk, R=>rst);
   lat_label_2_input_9 : latch port map ( Q=>label_2_input_9, D=>nx4702, CLK
      =>nx34549);
   reg_label_2_input_state_machine_9 : dffr port map ( Q=>
      label_2_input_state_machine_9, QB=>OPEN, D=>nx16543, CLK=>clk, R=>rst
   );
   ix4699 : xnor2 port map ( Y=>nx4698, A0=>nx4688, A1=>nx33443);
   ix4689 : oai22 port map ( Y=>nx4688, A0=>nx33338, A1=>nx33432, B0=>
      nx33442, B1=>nx28602);
   ix33339 : aoi22 port map ( Y=>nx33338, A0=>label_2_output(7), A1=>
      booth_booth_integration_output_1_7, B0=>nx4624, B1=>nx13051);
   labelsregfile_label2_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_2_output(7), QB=>OPEN, D=>nx16513, CLK=>clk, R=>rst);
   lat_label_2_input_7 : latch port map ( Q=>label_2_input_7, D=>nx4638, CLK
      =>nx34549);
   reg_label_2_input_state_machine_7 : dffr port map ( Q=>
      label_2_input_state_machine_7, QB=>OPEN, D=>nx16503, CLK=>clk, R=>rst
   );
   ix4635 : xnor2 port map ( Y=>nx4634, A0=>nx4624, A1=>nx33428);
   ix4625 : oai22 port map ( Y=>nx4624, A0=>nx33349, A1=>nx33417, B0=>
      nx33427, B1=>nx28604);
   ix33350 : aoi22 port map ( Y=>nx33349, A0=>label_2_output(5), A1=>
      booth_booth_integration_output_1_5, B0=>nx4560, B1=>nx13049);
   labelsregfile_label2_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_2_output(5), QB=>OPEN, D=>nx16473, CLK=>clk, R=>rst);
   lat_label_2_input_5 : latch port map ( Q=>label_2_input_5, D=>nx4574, CLK
      =>nx34549);
   reg_label_2_input_state_machine_5 : dffr port map ( Q=>
      label_2_input_state_machine_5, QB=>OPEN, D=>nx16463, CLK=>clk, R=>rst
   );
   ix4571 : xnor2 port map ( Y=>nx4570, A0=>nx4560, A1=>nx33413);
   ix4561 : oai22 port map ( Y=>nx4560, A0=>nx33360, A1=>nx33402, B0=>
      nx33412, B1=>nx28606);
   ix33361 : aoi22 port map ( Y=>nx33360, A0=>label_2_output(3), A1=>
      booth_booth_integration_output_1_3, B0=>nx4496, B1=>nx13045);
   labelsregfile_label2_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_2_output(3), QB=>OPEN, D=>nx16433, CLK=>clk, R=>rst);
   lat_label_2_input_3 : latch port map ( Q=>label_2_input_3, D=>nx4510, CLK
      =>nx34547);
   reg_label_2_input_state_machine_3 : dffr port map ( Q=>
      label_2_input_state_machine_3, QB=>OPEN, D=>nx16423, CLK=>clk, R=>rst
   );
   ix4507 : xnor2 port map ( Y=>nx4506, A0=>nx4496, A1=>nx33398);
   ix4497 : oai22 port map ( Y=>nx4496, A0=>nx33371, A1=>nx33387, B0=>
      nx33397, B1=>nx28608);
   ix33372 : aoi32 port map ( Y=>nx33371, A0=>label_2_output(0), A1=>nx35727, 
      A2=>nx13042, B0=>label_2_output(1), B1=>
      booth_booth_integration_output_1_1);
   labelsregfile_label2_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_2_output(1), QB=>OPEN, D=>nx16393, CLK=>clk, R=>rst);
   lat_label_2_input_1 : latch port map ( Q=>label_2_input_1, D=>nx4446, CLK
      =>nx34547);
   reg_label_2_input_state_machine_1 : dffr port map ( Q=>
      label_2_input_state_machine_1, QB=>OPEN, D=>nx16383, CLK=>clk, R=>rst
   );
   ix4443 : xor2 port map ( Y=>nx4442, A0=>nx33382, A1=>nx33384);
   ix33383 : nand02 port map ( Y=>nx33382, A0=>label_2_output(0), A1=>
      nx35727);
   ix33385 : xnor2 port map ( Y=>nx33384, A0=>
      booth_booth_integration_output_1_1, A1=>label_2_output(1));
   labelsregfile_label2_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_2_output(2), QB=>nx33397, D=>nx16413, CLK=>clk, R=>rst);
   lat_label_2_input_2 : latch port map ( Q=>label_2_input_2, D=>nx4478, CLK
      =>nx34547);
   reg_label_2_input_state_machine_2 : dffr port map ( Q=>
      label_2_input_state_machine_2, QB=>OPEN, D=>nx16403, CLK=>clk, R=>rst
   );
   ix4475 : xor2 port map ( Y=>nx4474, A0=>nx33371, A1=>nx33387);
   ix33399 : xnor2 port map ( Y=>nx33398, A0=>
      booth_booth_integration_output_1_3, A1=>label_2_output(3));
   labelsregfile_label2_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_2_output(4), QB=>nx33412, D=>nx16453, CLK=>clk, R=>rst);
   lat_label_2_input_4 : latch port map ( Q=>label_2_input_4, D=>nx4542, CLK
      =>nx34549);
   reg_label_2_input_state_machine_4 : dffr port map ( Q=>
      label_2_input_state_machine_4, QB=>OPEN, D=>nx16443, CLK=>clk, R=>rst
   );
   ix4539 : xor2 port map ( Y=>nx4538, A0=>nx33360, A1=>nx33402);
   ix33414 : xnor2 port map ( Y=>nx33413, A0=>
      booth_booth_integration_output_1_5, A1=>label_2_output(5));
   labelsregfile_label2_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_2_output(6), QB=>nx33427, D=>nx16493, CLK=>clk, R=>rst);
   lat_label_2_input_6 : latch port map ( Q=>label_2_input_6, D=>nx4606, CLK
      =>nx34549);
   reg_label_2_input_state_machine_6 : dffr port map ( Q=>
      label_2_input_state_machine_6, QB=>OPEN, D=>nx16483, CLK=>clk, R=>rst
   );
   ix4603 : xor2 port map ( Y=>nx4602, A0=>nx33349, A1=>nx33417);
   ix33429 : xnor2 port map ( Y=>nx33428, A0=>
      booth_booth_integration_output_1_7, A1=>label_2_output(7));
   labelsregfile_label2_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_2_output(8), QB=>nx33442, D=>nx16533, CLK=>clk, R=>rst);
   lat_label_2_input_8 : latch port map ( Q=>label_2_input_8, D=>nx4670, CLK
      =>nx34549);
   reg_label_2_input_state_machine_8 : dffr port map ( Q=>
      label_2_input_state_machine_8, QB=>OPEN, D=>nx16523, CLK=>clk, R=>rst
   );
   ix4667 : xor2 port map ( Y=>nx4666, A0=>nx33338, A1=>nx33432);
   ix33444 : xnor2 port map ( Y=>nx33443, A0=>
      booth_booth_integration_output_1_9, A1=>label_2_output(9));
   labelsregfile_label2_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_2_output(10), QB=>nx33457, D=>nx16573, CLK=>clk, R=>rst);
   lat_label_2_input_10 : latch port map ( Q=>label_2_input_10, D=>nx4734, 
      CLK=>nx34549);
   reg_label_2_input_state_machine_10 : dffr port map ( Q=>
      label_2_input_state_machine_10, QB=>OPEN, D=>nx16563, CLK=>clk, R=>rst
   );
   ix4731 : xor2 port map ( Y=>nx4730, A0=>nx33327, A1=>nx33447);
   ix33459 : xnor2 port map ( Y=>nx33458, A0=>
      booth_booth_integration_output_1_11, A1=>label_2_output(11));
   labelsregfile_label2_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_2_output(12), QB=>nx33472, D=>nx16613, CLK=>clk, R=>rst);
   lat_label_2_input_12 : latch port map ( Q=>label_2_input_12, D=>nx4798, 
      CLK=>nx34551);
   reg_label_2_input_state_machine_12 : dffr port map ( Q=>
      label_2_input_state_machine_12, QB=>OPEN, D=>nx16603, CLK=>clk, R=>rst
   );
   ix4795 : xor2 port map ( Y=>nx4794, A0=>nx33316, A1=>nx33462);
   ix33474 : xnor2 port map ( Y=>nx33473, A0=>
      booth_booth_integration_output_1_13, A1=>label_2_output(13));
   max_calc_reg_ans2_14 : dff port map ( Q=>max_calc_ans2_14, QB=>OPEN, D=>
      nx24323, CLK=>clk);
   max_calc_reg_ans7_14 : dff port map ( Q=>max_calc_ans7_14, QB=>OPEN, D=>
      nx24383, CLK=>clk);
   max_calc_reg_ans8_14 : dff port map ( Q=>max_calc_ans8_14, QB=>OPEN, D=>
      nx24373, CLK=>clk);
   max_calc_reg_comparator_first_inp1_14 : dff port map ( Q=>
      max_calc_comparator_first_inp1_14, QB=>OPEN, D=>nx24363, CLK=>clk);
   labelsregfile_label1_loop1_14_fx_reg_q : dffr port map ( Q=>
      label_1_output(14), QB=>nx33677, D=>nx17503, CLK=>clk, R=>rst);
   lat_label_1_input_14 : latch port map ( Q=>label_1_input_14, D=>nx6200, 
      CLK=>nx34555);
   reg_label_1_input_state_machine_14 : dffr port map ( Q=>
      label_1_input_state_machine_14, QB=>OPEN, D=>nx17493, CLK=>clk, R=>rst
   );
   ix6197 : xor2 port map ( Y=>nx6196, A0=>nx33503, A1=>nx33675);
   ix33504 : aoi22 port map ( Y=>nx33503, A0=>label_1_output(13), A1=>
      booth_booth_integration_output_0_13, B0=>nx6154, B1=>nx13114);
   labelsregfile_label1_loop1_13_fx_reg_q : dffr port map ( Q=>
      label_1_output(13), QB=>OPEN, D=>nx17483, CLK=>clk, R=>rst);
   lat_label_1_input_13 : latch port map ( Q=>label_1_input_13, D=>nx6168, 
      CLK=>nx34555);
   reg_label_1_input_state_machine_13 : dffr port map ( Q=>
      label_1_input_state_machine_13, QB=>OPEN, D=>nx17473, CLK=>clk, R=>rst
   );
   ix6165 : xnor2 port map ( Y=>nx6164, A0=>nx6154, A1=>nx33671);
   ix6155 : oai22 port map ( Y=>nx6154, A0=>nx33514, A1=>nx33660, B0=>
      nx33670, B1=>nx26638);
   ix33515 : aoi22 port map ( Y=>nx33514, A0=>label_1_output(11), A1=>
      booth_booth_integration_output_0_11, B0=>nx6090, B1=>nx13111);
   labelsregfile_label1_loop1_11_fx_reg_q : dffr port map ( Q=>
      label_1_output(11), QB=>OPEN, D=>nx17443, CLK=>clk, R=>rst);
   lat_label_1_input_11 : latch port map ( Q=>label_1_input_11, D=>nx6104, 
      CLK=>nx34555);
   reg_label_1_input_state_machine_11 : dffr port map ( Q=>
      label_1_input_state_machine_11, QB=>OPEN, D=>nx17433, CLK=>clk, R=>rst
   );
   ix6101 : xnor2 port map ( Y=>nx6100, A0=>nx6090, A1=>nx33656);
   ix6091 : oai22 port map ( Y=>nx6090, A0=>nx33525, A1=>nx33645, B0=>
      nx33655, B1=>nx26640);
   ix33526 : aoi22 port map ( Y=>nx33525, A0=>label_1_output(9), A1=>
      booth_booth_integration_output_0_9, B0=>nx6026, B1=>nx13107);
   labelsregfile_label1_loop1_9_fx_reg_q : dffr port map ( Q=>
      label_1_output(9), QB=>OPEN, D=>nx17403, CLK=>clk, R=>rst);
   lat_label_1_input_9 : latch port map ( Q=>label_1_input_9, D=>nx6040, CLK
      =>nx34553);
   reg_label_1_input_state_machine_9 : dffr port map ( Q=>
      label_1_input_state_machine_9, QB=>OPEN, D=>nx17393, CLK=>clk, R=>rst
   );
   ix6037 : xnor2 port map ( Y=>nx6036, A0=>nx6026, A1=>nx33641);
   ix6027 : oai22 port map ( Y=>nx6026, A0=>nx33536, A1=>nx33630, B0=>
      nx33640, B1=>nx26642);
   ix33537 : aoi22 port map ( Y=>nx33536, A0=>label_1_output(7), A1=>
      booth_booth_integration_output_0_7, B0=>nx5962, B1=>nx13103);
   labelsregfile_label1_loop1_7_fx_reg_q : dffr port map ( Q=>
      label_1_output(7), QB=>OPEN, D=>nx17363, CLK=>clk, R=>rst);
   lat_label_1_input_7 : latch port map ( Q=>label_1_input_7, D=>nx5976, CLK
      =>nx34553);
   reg_label_1_input_state_machine_7 : dffr port map ( Q=>
      label_1_input_state_machine_7, QB=>OPEN, D=>nx17353, CLK=>clk, R=>rst
   );
   ix5973 : xnor2 port map ( Y=>nx5972, A0=>nx5962, A1=>nx33626);
   ix5963 : oai22 port map ( Y=>nx5962, A0=>nx33547, A1=>nx33615, B0=>
      nx33625, B1=>nx26644);
   ix33548 : aoi22 port map ( Y=>nx33547, A0=>label_1_output(5), A1=>
      booth_booth_integration_output_0_5, B0=>nx5898, B1=>nx13099);
   labelsregfile_label1_loop1_5_fx_reg_q : dffr port map ( Q=>
      label_1_output(5), QB=>OPEN, D=>nx17323, CLK=>clk, R=>rst);
   lat_label_1_input_5 : latch port map ( Q=>label_1_input_5, D=>nx5912, CLK
      =>nx34553);
   reg_label_1_input_state_machine_5 : dffr port map ( Q=>
      label_1_input_state_machine_5, QB=>OPEN, D=>nx17313, CLK=>clk, R=>rst
   );
   ix5909 : xnor2 port map ( Y=>nx5908, A0=>nx5898, A1=>nx33611);
   ix5899 : oai22 port map ( Y=>nx5898, A0=>nx33558, A1=>nx33600, B0=>
      nx33610, B1=>nx26646);
   ix33559 : aoi22 port map ( Y=>nx33558, A0=>label_1_output(3), A1=>
      booth_booth_integration_output_0_3, B0=>nx5834, B1=>nx13097);
   labelsregfile_label1_loop1_3_fx_reg_q : dffr port map ( Q=>
      label_1_output(3), QB=>OPEN, D=>nx17283, CLK=>clk, R=>rst);
   lat_label_1_input_3 : latch port map ( Q=>label_1_input_3, D=>nx5848, CLK
      =>nx34551);
   reg_label_1_input_state_machine_3 : dffr port map ( Q=>
      label_1_input_state_machine_3, QB=>OPEN, D=>nx17273, CLK=>clk, R=>rst
   );
   ix5845 : xnor2 port map ( Y=>nx5844, A0=>nx5834, A1=>nx33596);
   ix5835 : oai22 port map ( Y=>nx5834, A0=>nx33569, A1=>nx33585, B0=>
      nx33595, B1=>nx26648);
   ix33570 : aoi32 port map ( Y=>nx33569, A0=>label_1_output(0), A1=>nx35731, 
      A2=>nx13093, B0=>label_1_output(1), B1=>
      booth_booth_integration_output_0_1);
   labelsregfile_label1_loop1_1_fx_reg_q : dffr port map ( Q=>
      label_1_output(1), QB=>OPEN, D=>nx17243, CLK=>clk, R=>rst);
   lat_label_1_input_1 : latch port map ( Q=>label_1_input_1, D=>nx5784, CLK
      =>nx34551);
   reg_label_1_input_state_machine_1 : dffr port map ( Q=>
      label_1_input_state_machine_1, QB=>OPEN, D=>nx17233, CLK=>clk, R=>rst
   );
   ix5781 : xor2 port map ( Y=>nx5780, A0=>nx33580, A1=>nx33582);
   ix33581 : nand02 port map ( Y=>nx33580, A0=>label_1_output(0), A1=>
      nx35731);
   ix33583 : xnor2 port map ( Y=>nx33582, A0=>
      booth_booth_integration_output_0_1, A1=>label_1_output(1));
   labelsregfile_label1_loop1_2_fx_reg_q : dffr port map ( Q=>
      label_1_output(2), QB=>nx33595, D=>nx17263, CLK=>clk, R=>rst);
   lat_label_1_input_2 : latch port map ( Q=>label_1_input_2, D=>nx5816, CLK
      =>nx34551);
   reg_label_1_input_state_machine_2 : dffr port map ( Q=>
      label_1_input_state_machine_2, QB=>OPEN, D=>nx17253, CLK=>clk, R=>rst
   );
   ix5813 : xor2 port map ( Y=>nx5812, A0=>nx33569, A1=>nx33585);
   ix33597 : xnor2 port map ( Y=>nx33596, A0=>
      booth_booth_integration_output_0_3, A1=>label_1_output(3));
   labelsregfile_label1_loop1_4_fx_reg_q : dffr port map ( Q=>
      label_1_output(4), QB=>nx33610, D=>nx17303, CLK=>clk, R=>rst);
   lat_label_1_input_4 : latch port map ( Q=>label_1_input_4, D=>nx5880, CLK
      =>nx34553);
   reg_label_1_input_state_machine_4 : dffr port map ( Q=>
      label_1_input_state_machine_4, QB=>OPEN, D=>nx17293, CLK=>clk, R=>rst
   );
   ix5877 : xor2 port map ( Y=>nx5876, A0=>nx33558, A1=>nx33600);
   ix33612 : xnor2 port map ( Y=>nx33611, A0=>
      booth_booth_integration_output_0_5, A1=>label_1_output(5));
   labelsregfile_label1_loop1_6_fx_reg_q : dffr port map ( Q=>
      label_1_output(6), QB=>nx33625, D=>nx17343, CLK=>clk, R=>rst);
   lat_label_1_input_6 : latch port map ( Q=>label_1_input_6, D=>nx5944, CLK
      =>nx34553);
   reg_label_1_input_state_machine_6 : dffr port map ( Q=>
      label_1_input_state_machine_6, QB=>OPEN, D=>nx17333, CLK=>clk, R=>rst
   );
   ix5941 : xor2 port map ( Y=>nx5940, A0=>nx33547, A1=>nx33615);
   ix33627 : xnor2 port map ( Y=>nx33626, A0=>
      booth_booth_integration_output_0_7, A1=>label_1_output(7));
   labelsregfile_label1_loop1_8_fx_reg_q : dffr port map ( Q=>
      label_1_output(8), QB=>nx33640, D=>nx17383, CLK=>clk, R=>rst);
   lat_label_1_input_8 : latch port map ( Q=>label_1_input_8, D=>nx6008, CLK
      =>nx34553);
   reg_label_1_input_state_machine_8 : dffr port map ( Q=>
      label_1_input_state_machine_8, QB=>OPEN, D=>nx17373, CLK=>clk, R=>rst
   );
   ix6005 : xor2 port map ( Y=>nx6004, A0=>nx33536, A1=>nx33630);
   ix33642 : xnor2 port map ( Y=>nx33641, A0=>
      booth_booth_integration_output_0_9, A1=>label_1_output(9));
   labelsregfile_label1_loop1_10_fx_reg_q : dffr port map ( Q=>
      label_1_output(10), QB=>nx33655, D=>nx17423, CLK=>clk, R=>rst);
   lat_label_1_input_10 : latch port map ( Q=>label_1_input_10, D=>nx6072, 
      CLK=>nx34553);
   reg_label_1_input_state_machine_10 : dffr port map ( Q=>
      label_1_input_state_machine_10, QB=>OPEN, D=>nx17413, CLK=>clk, R=>rst
   );
   ix6069 : xor2 port map ( Y=>nx6068, A0=>nx33525, A1=>nx33645);
   ix33657 : xnor2 port map ( Y=>nx33656, A0=>
      booth_booth_integration_output_0_11, A1=>label_1_output(11));
   labelsregfile_label1_loop1_12_fx_reg_q : dffr port map ( Q=>
      label_1_output(12), QB=>nx33670, D=>nx17463, CLK=>clk, R=>rst);
   lat_label_1_input_12 : latch port map ( Q=>label_1_input_12, D=>nx6136, 
      CLK=>nx34555);
   reg_label_1_input_state_machine_12 : dffr port map ( Q=>
      label_1_input_state_machine_12, QB=>OPEN, D=>nx17453, CLK=>clk, R=>rst
   );
   ix6133 : xor2 port map ( Y=>nx6132, A0=>nx33514, A1=>nx33660);
   ix33672 : xnor2 port map ( Y=>nx33671, A0=>
      booth_booth_integration_output_0_13, A1=>label_1_output(13));
   max_calc_reg_ans1_14 : dff port map ( Q=>max_calc_ans1_14, QB=>OPEN, D=>
      nx24333, CLK=>clk);
   max_calc_reg_ans6_14 : dff port map ( Q=>max_calc_ans6_14, QB=>OPEN, D=>
      nx24343, CLK=>clk);
   max_calc_reg_ans5_14 : dff port map ( Q=>max_calc_ans5_14, QB=>OPEN, D=>
      nx24353, CLK=>clk);
   max_calc_reg_comparator_first_inp2_14 : dff port map ( Q=>
      max_calc_comparator_first_inp2_14, QB=>nx33292, D=>nx24393, CLK=>clk);
   ix19011 : oai22 port map ( Y=>nx19010, A0=>nx33694, A1=>nx33729, B0=>
      max_calc_comparator_first_inp2_13, B1=>nx33726);
   max_calc_reg_comparator_first_inp2_13 : dff port map ( Q=>
      max_calc_comparator_first_inp2_13, QB=>OPEN, D=>nx24473, CLK=>clk);
   max_calc_reg_ans2_13 : dff port map ( Q=>max_calc_ans2_13, QB=>OPEN, D=>
      nx24403, CLK=>clk);
   max_calc_reg_ans7_13 : dff port map ( Q=>max_calc_ans7_13, QB=>OPEN, D=>
      nx24463, CLK=>clk);
   max_calc_reg_ans8_13 : dff port map ( Q=>max_calc_ans8_13, QB=>OPEN, D=>
      nx24453, CLK=>clk);
   max_calc_reg_comparator_first_inp1_13 : dff port map ( Q=>
      max_calc_comparator_first_inp1_13, QB=>nx33726, D=>nx24443, CLK=>clk);
   max_calc_reg_ans1_13 : dff port map ( Q=>max_calc_ans1_13, QB=>OPEN, D=>
      nx24413, CLK=>clk);
   max_calc_reg_ans6_13 : dff port map ( Q=>max_calc_ans6_13, QB=>OPEN, D=>
      nx24423, CLK=>clk);
   max_calc_reg_ans5_13 : dff port map ( Q=>max_calc_ans5_13, QB=>OPEN, D=>
      nx24433, CLK=>clk);
   ix33730 : aoi22 port map ( Y=>nx33729, A0=>nx33731, A1=>
      max_calc_comparator_first_inp1_12, B0=>nx17500, B1=>nx18994);
   max_calc_reg_ans2_12 : dff port map ( Q=>max_calc_ans2_12, QB=>OPEN, D=>
      nx24483, CLK=>clk);
   max_calc_reg_ans7_12 : dff port map ( Q=>max_calc_ans7_12, QB=>OPEN, D=>
      nx24543, CLK=>clk);
   max_calc_reg_ans8_12 : dff port map ( Q=>max_calc_ans8_12, QB=>OPEN, D=>
      nx24533, CLK=>clk);
   max_calc_reg_comparator_first_inp1_12 : dff port map ( Q=>
      max_calc_comparator_first_inp1_12, QB=>OPEN, D=>nx24523, CLK=>clk);
   max_calc_reg_ans1_12 : dff port map ( Q=>max_calc_ans1_12, QB=>OPEN, D=>
      nx24493, CLK=>clk);
   max_calc_reg_ans6_12 : dff port map ( Q=>max_calc_ans6_12, QB=>OPEN, D=>
      nx24503, CLK=>clk);
   max_calc_reg_ans5_12 : dff port map ( Q=>max_calc_ans5_12, QB=>OPEN, D=>
      nx24513, CLK=>clk);
   max_calc_reg_comparator_first_inp2_12 : dff port map ( Q=>
      max_calc_comparator_first_inp2_12, QB=>nx33731, D=>nx24553, CLK=>clk);
   ix18995 : oai22 port map ( Y=>nx18994, A0=>nx33767, A1=>nx33802, B0=>
      max_calc_comparator_first_inp2_11, B1=>nx33799);
   max_calc_reg_comparator_first_inp2_11 : dff port map ( Q=>
      max_calc_comparator_first_inp2_11, QB=>OPEN, D=>nx24633, CLK=>clk);
   max_calc_reg_ans2_11 : dff port map ( Q=>max_calc_ans2_11, QB=>OPEN, D=>
      nx24563, CLK=>clk);
   max_calc_reg_ans7_11 : dff port map ( Q=>max_calc_ans7_11, QB=>OPEN, D=>
      nx24623, CLK=>clk);
   max_calc_reg_ans8_11 : dff port map ( Q=>max_calc_ans8_11, QB=>OPEN, D=>
      nx24613, CLK=>clk);
   max_calc_reg_comparator_first_inp1_11 : dff port map ( Q=>
      max_calc_comparator_first_inp1_11, QB=>nx33799, D=>nx24603, CLK=>clk);
   max_calc_reg_ans1_11 : dff port map ( Q=>max_calc_ans1_11, QB=>OPEN, D=>
      nx24573, CLK=>clk);
   max_calc_reg_ans6_11 : dff port map ( Q=>max_calc_ans6_11, QB=>OPEN, D=>
      nx24583, CLK=>clk);
   max_calc_reg_ans5_11 : dff port map ( Q=>max_calc_ans5_11, QB=>OPEN, D=>
      nx24593, CLK=>clk);
   ix33803 : aoi22 port map ( Y=>nx33802, A0=>nx33804, A1=>
      max_calc_comparator_first_inp1_10, B0=>nx17744, B1=>nx18978);
   max_calc_reg_ans2_10 : dff port map ( Q=>max_calc_ans2_10, QB=>OPEN, D=>
      nx24643, CLK=>clk);
   max_calc_reg_ans7_10 : dff port map ( Q=>max_calc_ans7_10, QB=>OPEN, D=>
      nx24703, CLK=>clk);
   max_calc_reg_ans8_10 : dff port map ( Q=>max_calc_ans8_10, QB=>OPEN, D=>
      nx24693, CLK=>clk);
   max_calc_reg_comparator_first_inp1_10 : dff port map ( Q=>
      max_calc_comparator_first_inp1_10, QB=>OPEN, D=>nx24683, CLK=>clk);
   max_calc_reg_ans1_10 : dff port map ( Q=>max_calc_ans1_10, QB=>OPEN, D=>
      nx24653, CLK=>clk);
   max_calc_reg_ans6_10 : dff port map ( Q=>max_calc_ans6_10, QB=>OPEN, D=>
      nx24663, CLK=>clk);
   max_calc_reg_ans5_10 : dff port map ( Q=>max_calc_ans5_10, QB=>OPEN, D=>
      nx24673, CLK=>clk);
   max_calc_reg_comparator_first_inp2_10 : dff port map ( Q=>
      max_calc_comparator_first_inp2_10, QB=>nx33804, D=>nx24713, CLK=>clk);
   ix18979 : oai22 port map ( Y=>nx18978, A0=>nx33840, A1=>nx33875, B0=>
      max_calc_comparator_first_inp2_9, B1=>nx33872);
   max_calc_reg_comparator_first_inp2_9 : dff port map ( Q=>
      max_calc_comparator_first_inp2_9, QB=>OPEN, D=>nx24793, CLK=>clk);
   max_calc_reg_ans2_9 : dff port map ( Q=>max_calc_ans2_9, QB=>OPEN, D=>
      nx24723, CLK=>clk);
   max_calc_reg_ans7_9 : dff port map ( Q=>max_calc_ans7_9, QB=>OPEN, D=>
      nx24783, CLK=>clk);
   max_calc_reg_ans8_9 : dff port map ( Q=>max_calc_ans8_9, QB=>OPEN, D=>
      nx24773, CLK=>clk);
   max_calc_reg_comparator_first_inp1_9 : dff port map ( Q=>
      max_calc_comparator_first_inp1_9, QB=>nx33872, D=>nx24763, CLK=>clk);
   max_calc_reg_ans1_9 : dff port map ( Q=>max_calc_ans1_9, QB=>OPEN, D=>
      nx24733, CLK=>clk);
   max_calc_reg_ans6_9 : dff port map ( Q=>max_calc_ans6_9, QB=>OPEN, D=>
      nx24743, CLK=>clk);
   max_calc_reg_ans5_9 : dff port map ( Q=>max_calc_ans5_9, QB=>OPEN, D=>
      nx24753, CLK=>clk);
   ix33876 : aoi22 port map ( Y=>nx33875, A0=>nx33877, A1=>
      max_calc_comparator_first_inp1_8, B0=>nx17988, B1=>nx18962);
   max_calc_reg_ans2_8 : dff port map ( Q=>max_calc_ans2_8, QB=>OPEN, D=>
      nx24803, CLK=>clk);
   max_calc_reg_ans7_8 : dff port map ( Q=>max_calc_ans7_8, QB=>OPEN, D=>
      nx24863, CLK=>clk);
   max_calc_reg_ans8_8 : dff port map ( Q=>max_calc_ans8_8, QB=>OPEN, D=>
      nx24853, CLK=>clk);
   max_calc_reg_comparator_first_inp1_8 : dff port map ( Q=>
      max_calc_comparator_first_inp1_8, QB=>OPEN, D=>nx24843, CLK=>clk);
   max_calc_reg_ans1_8 : dff port map ( Q=>max_calc_ans1_8, QB=>OPEN, D=>
      nx24813, CLK=>clk);
   max_calc_reg_ans6_8 : dff port map ( Q=>max_calc_ans6_8, QB=>OPEN, D=>
      nx24823, CLK=>clk);
   max_calc_reg_ans5_8 : dff port map ( Q=>max_calc_ans5_8, QB=>OPEN, D=>
      nx24833, CLK=>clk);
   max_calc_reg_comparator_first_inp2_8 : dff port map ( Q=>
      max_calc_comparator_first_inp2_8, QB=>nx33877, D=>nx24873, CLK=>clk);
   ix18963 : oai22 port map ( Y=>nx18962, A0=>nx33913, A1=>nx33948, B0=>
      max_calc_comparator_first_inp2_7, B1=>nx33945);
   max_calc_reg_comparator_first_inp2_7 : dff port map ( Q=>
      max_calc_comparator_first_inp2_7, QB=>OPEN, D=>nx24953, CLK=>clk);
   max_calc_reg_ans2_7 : dff port map ( Q=>max_calc_ans2_7, QB=>OPEN, D=>
      nx24883, CLK=>clk);
   max_calc_reg_ans7_7 : dff port map ( Q=>max_calc_ans7_7, QB=>OPEN, D=>
      nx24943, CLK=>clk);
   max_calc_reg_ans8_7 : dff port map ( Q=>max_calc_ans8_7, QB=>OPEN, D=>
      nx24933, CLK=>clk);
   max_calc_reg_comparator_first_inp1_7 : dff port map ( Q=>
      max_calc_comparator_first_inp1_7, QB=>nx33945, D=>nx24923, CLK=>clk);
   max_calc_reg_ans1_7 : dff port map ( Q=>max_calc_ans1_7, QB=>OPEN, D=>
      nx24893, CLK=>clk);
   max_calc_reg_ans6_7 : dff port map ( Q=>max_calc_ans6_7, QB=>OPEN, D=>
      nx24903, CLK=>clk);
   max_calc_reg_ans5_7 : dff port map ( Q=>max_calc_ans5_7, QB=>OPEN, D=>
      nx24913, CLK=>clk);
   ix33949 : aoi22 port map ( Y=>nx33948, A0=>nx33950, A1=>
      max_calc_comparator_first_inp1_6, B0=>nx18232, B1=>nx18946);
   max_calc_reg_ans2_6 : dff port map ( Q=>max_calc_ans2_6, QB=>OPEN, D=>
      nx24963, CLK=>clk);
   max_calc_reg_ans7_6 : dff port map ( Q=>max_calc_ans7_6, QB=>OPEN, D=>
      nx25023, CLK=>clk);
   max_calc_reg_ans8_6 : dff port map ( Q=>max_calc_ans8_6, QB=>OPEN, D=>
      nx25013, CLK=>clk);
   max_calc_reg_comparator_first_inp1_6 : dff port map ( Q=>
      max_calc_comparator_first_inp1_6, QB=>OPEN, D=>nx25003, CLK=>clk);
   max_calc_reg_ans1_6 : dff port map ( Q=>max_calc_ans1_6, QB=>OPEN, D=>
      nx24973, CLK=>clk);
   max_calc_reg_ans6_6 : dff port map ( Q=>max_calc_ans6_6, QB=>OPEN, D=>
      nx24983, CLK=>clk);
   max_calc_reg_ans5_6 : dff port map ( Q=>max_calc_ans5_6, QB=>OPEN, D=>
      nx24993, CLK=>clk);
   max_calc_reg_comparator_first_inp2_6 : dff port map ( Q=>
      max_calc_comparator_first_inp2_6, QB=>nx33950, D=>nx25033, CLK=>clk);
   ix18947 : oai22 port map ( Y=>nx18946, A0=>nx33986, A1=>nx34021, B0=>
      max_calc_comparator_first_inp2_5, B1=>nx34018);
   max_calc_reg_comparator_first_inp2_5 : dff port map ( Q=>
      max_calc_comparator_first_inp2_5, QB=>OPEN, D=>nx25113, CLK=>clk);
   max_calc_reg_ans2_5 : dff port map ( Q=>max_calc_ans2_5, QB=>OPEN, D=>
      nx25043, CLK=>clk);
   max_calc_reg_ans7_5 : dff port map ( Q=>max_calc_ans7_5, QB=>OPEN, D=>
      nx25103, CLK=>clk);
   max_calc_reg_ans8_5 : dff port map ( Q=>max_calc_ans8_5, QB=>OPEN, D=>
      nx25093, CLK=>clk);
   max_calc_reg_comparator_first_inp1_5 : dff port map ( Q=>
      max_calc_comparator_first_inp1_5, QB=>nx34018, D=>nx25083, CLK=>clk);
   max_calc_reg_ans1_5 : dff port map ( Q=>max_calc_ans1_5, QB=>OPEN, D=>
      nx25053, CLK=>clk);
   max_calc_reg_ans6_5 : dff port map ( Q=>max_calc_ans6_5, QB=>OPEN, D=>
      nx25063, CLK=>clk);
   max_calc_reg_ans5_5 : dff port map ( Q=>max_calc_ans5_5, QB=>OPEN, D=>
      nx25073, CLK=>clk);
   ix34022 : aoi22 port map ( Y=>nx34021, A0=>nx34023, A1=>
      max_calc_comparator_first_inp1_4, B0=>nx18476, B1=>nx18930);
   max_calc_reg_ans2_4 : dff port map ( Q=>max_calc_ans2_4, QB=>OPEN, D=>
      nx25123, CLK=>clk);
   max_calc_reg_ans7_4 : dff port map ( Q=>max_calc_ans7_4, QB=>OPEN, D=>
      nx25183, CLK=>clk);
   max_calc_reg_ans8_4 : dff port map ( Q=>max_calc_ans8_4, QB=>OPEN, D=>
      nx25173, CLK=>clk);
   max_calc_reg_comparator_first_inp1_4 : dff port map ( Q=>
      max_calc_comparator_first_inp1_4, QB=>OPEN, D=>nx25163, CLK=>clk);
   max_calc_reg_ans1_4 : dff port map ( Q=>max_calc_ans1_4, QB=>OPEN, D=>
      nx25133, CLK=>clk);
   max_calc_reg_ans6_4 : dff port map ( Q=>max_calc_ans6_4, QB=>OPEN, D=>
      nx25143, CLK=>clk);
   max_calc_reg_ans5_4 : dff port map ( Q=>max_calc_ans5_4, QB=>OPEN, D=>
      nx25153, CLK=>clk);
   max_calc_reg_comparator_first_inp2_4 : dff port map ( Q=>
      max_calc_comparator_first_inp2_4, QB=>nx34023, D=>nx25193, CLK=>clk);
   ix18931 : oai22 port map ( Y=>nx18930, A0=>nx34059, A1=>nx34094, B0=>
      max_calc_comparator_first_inp2_3, B1=>nx34091);
   max_calc_reg_comparator_first_inp2_3 : dff port map ( Q=>
      max_calc_comparator_first_inp2_3, QB=>OPEN, D=>nx25273, CLK=>clk);
   max_calc_reg_ans2_3 : dff port map ( Q=>max_calc_ans2_3, QB=>OPEN, D=>
      nx25203, CLK=>clk);
   max_calc_reg_ans7_3 : dff port map ( Q=>max_calc_ans7_3, QB=>OPEN, D=>
      nx25263, CLK=>clk);
   max_calc_reg_ans8_3 : dff port map ( Q=>max_calc_ans8_3, QB=>OPEN, D=>
      nx25253, CLK=>clk);
   max_calc_reg_comparator_first_inp1_3 : dff port map ( Q=>
      max_calc_comparator_first_inp1_3, QB=>nx34091, D=>nx25243, CLK=>clk);
   max_calc_reg_ans1_3 : dff port map ( Q=>max_calc_ans1_3, QB=>OPEN, D=>
      nx25213, CLK=>clk);
   max_calc_reg_ans6_3 : dff port map ( Q=>max_calc_ans6_3, QB=>OPEN, D=>
      nx25223, CLK=>clk);
   max_calc_reg_ans5_3 : dff port map ( Q=>max_calc_ans5_3, QB=>OPEN, D=>
      nx25233, CLK=>clk);
   ix34095 : aoi22 port map ( Y=>nx34094, A0=>nx34096, A1=>
      max_calc_comparator_first_inp1_2, B0=>nx18720, B1=>nx18914);
   max_calc_reg_ans2_2 : dff port map ( Q=>max_calc_ans2_2, QB=>OPEN, D=>
      nx25283, CLK=>clk);
   max_calc_reg_ans7_2 : dff port map ( Q=>max_calc_ans7_2, QB=>OPEN, D=>
      nx25343, CLK=>clk);
   max_calc_reg_ans8_2 : dff port map ( Q=>max_calc_ans8_2, QB=>OPEN, D=>
      nx25333, CLK=>clk);
   max_calc_reg_comparator_first_inp1_2 : dff port map ( Q=>
      max_calc_comparator_first_inp1_2, QB=>OPEN, D=>nx25323, CLK=>clk);
   max_calc_reg_ans1_2 : dff port map ( Q=>max_calc_ans1_2, QB=>OPEN, D=>
      nx25293, CLK=>clk);
   max_calc_reg_ans6_2 : dff port map ( Q=>max_calc_ans6_2, QB=>OPEN, D=>
      nx25303, CLK=>clk);
   max_calc_reg_ans5_2 : dff port map ( Q=>max_calc_ans5_2, QB=>OPEN, D=>
      nx25313, CLK=>clk);
   max_calc_reg_comparator_first_inp2_2 : dff port map ( Q=>
      max_calc_comparator_first_inp2_2, QB=>nx34096, D=>nx25353, CLK=>clk);
   ix18915 : oai21 port map ( Y=>nx18914, A0=>
      max_calc_comparator_first_inp2_1, A1=>nx34162, B0=>nx34165);
   max_calc_reg_comparator_first_inp2_1 : dff port map ( Q=>
      max_calc_comparator_first_inp2_1, QB=>OPEN, D=>nx25433, CLK=>clk);
   max_calc_reg_ans2_1 : dff port map ( Q=>max_calc_ans2_1, QB=>OPEN, D=>
      nx25363, CLK=>clk);
   max_calc_reg_ans7_1 : dff port map ( Q=>max_calc_ans7_1, QB=>OPEN, D=>
      nx25423, CLK=>clk);
   max_calc_reg_ans8_1 : dff port map ( Q=>max_calc_ans8_1, QB=>OPEN, D=>
      nx25413, CLK=>clk);
   max_calc_reg_comparator_first_inp1_1 : dff port map ( Q=>
      max_calc_comparator_first_inp1_1, QB=>nx34162, D=>nx25403, CLK=>clk);
   max_calc_reg_ans1_1 : dff port map ( Q=>max_calc_ans1_1, QB=>OPEN, D=>
      nx25373, CLK=>clk);
   max_calc_reg_ans6_1 : dff port map ( Q=>max_calc_ans6_1, QB=>OPEN, D=>
      nx25383, CLK=>clk);
   max_calc_reg_ans5_1 : dff port map ( Q=>max_calc_ans5_1, QB=>OPEN, D=>
      nx25393, CLK=>clk);
   ix34166 : oai21 port map ( Y=>nx34165, A0=>nx33288, A1=>
      max_calc_comparator_first_inp1_0, B0=>nx18842);
   ix19141 : xnor2 port map ( Y=>nx19140, A0=>
      max_calc_comparator_first_inp2_15, A1=>
      max_calc_comparator_first_inp1_15);
   max_calc_reg_comparator_first_inp2_15 : dff port map ( Q=>
      max_calc_comparator_first_inp2_15, QB=>OPEN, D=>nx25553, CLK=>clk);
   labelsregfile_label2_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_2_output(15), QB=>OPEN, D=>nx16663, CLK=>clk, R=>rst);
   lat_label_2_input_15 : latch port map ( Q=>label_2_input_15, D=>nx4888, 
      CLK=>nx34555);
   reg_label_2_input_state_machine_15 : dffr port map ( Q=>
      label_2_input_state_machine_15, QB=>OPEN, D=>nx15823, CLK=>clk, R=>rst
   );
   ix4885 : xnor2 port map ( Y=>nx4884, A0=>nx4880, A1=>nx34182);
   ix4881 : oai22 port map ( Y=>nx4880, A0=>nx33305, A1=>nx33477, B0=>
      nx33479, B1=>nx28596);
   max_calc_reg_ans2_15 : dff port map ( Q=>max_calc_ans2_15, QB=>OPEN, D=>
      nx25483, CLK=>clk);
   max_calc_reg_ans7_15 : dff port map ( Q=>max_calc_ans7_15, QB=>OPEN, D=>
      nx25543, CLK=>clk);
   max_calc_reg_ans8_15 : dff port map ( Q=>max_calc_ans8_15, QB=>OPEN, D=>
      nx25533, CLK=>clk);
   max_calc_reg_comparator_first_inp1_15 : dff port map ( Q=>
      max_calc_comparator_first_inp1_15, QB=>OPEN, D=>nx25523, CLK=>clk);
   labelsregfile_label1_loop1_15_fx_reg_q : dffr port map ( Q=>
      label_1_output(15), QB=>OPEN, D=>nx17513, CLK=>clk, R=>rst);
   lat_label_1_input_15 : latch port map ( Q=>label_1_input_15, D=>nx6226, 
      CLK=>nx34555);
   reg_label_1_input_state_machine_15 : dffr port map ( Q=>
      label_1_input_state_machine_15, QB=>OPEN, D=>nx16673, CLK=>clk, R=>rst
   );
   ix6223 : xnor2 port map ( Y=>nx6222, A0=>nx6218, A1=>nx34209);
   ix6219 : oai22 port map ( Y=>nx6218, A0=>nx33503, A1=>nx33675, B0=>
      nx33677, B1=>nx26636);
   max_calc_reg_ans1_15 : dff port map ( Q=>max_calc_ans1_15, QB=>OPEN, D=>
      nx25493, CLK=>clk);
   max_calc_reg_ans6_15 : dff port map ( Q=>max_calc_ans6_15, QB=>OPEN, D=>
      nx25503, CLK=>clk);
   max_calc_reg_ans5_15 : dff port map ( Q=>max_calc_ans5_15, QB=>OPEN, D=>
      nx25513, CLK=>clk);
   max_calc_reg_answer_1 : dffr port map ( Q=>answer_1_EXMPLR, QB=>OPEN, D=>
      nx25573, CLK=>clk, R=>rst);
   max_calc_reg_answer_2 : dffr port map ( Q=>answer_2_EXMPLR, QB=>OPEN, D=>
      nx25583, CLK=>clk, R=>rst);
   max_calc_reg_answer_3 : dffr port map ( Q=>answer_3_EXMPLR, QB=>OPEN, D=>
      nx25593, CLK=>clk, R=>rst);
   max_calc_reg_answer_4 : dffr port map ( Q=>answer_4_EXMPLR, QB=>OPEN, D=>
      nx25603, CLK=>clk, R=>rst);
   max_calc_reg_answer_5 : dffr port map ( Q=>answer_5_EXMPLR, QB=>OPEN, D=>
      nx25613, CLK=>clk, R=>rst);
   max_calc_reg_answer_6 : dffr port map ( Q=>answer_6_EXMPLR, QB=>OPEN, D=>
      nx25623, CLK=>clk, R=>rst);
   max_calc_reg_answer_7 : dffr port map ( Q=>answer_7_EXMPLR, QB=>OPEN, D=>
      nx25633, CLK=>clk, R=>rst);
   max_calc_reg_answer_8 : dffr port map ( Q=>answer_8_EXMPLR, QB=>OPEN, D=>
      nx25643, CLK=>clk, R=>rst);
   max_calc_reg_answer_9 : dffr port map ( Q=>answer_9_EXMPLR, QB=>OPEN, D=>
      nx25653, CLK=>clk, R=>rst);
   max_calc_reg_answer_10 : dffr port map ( Q=>answer_10_EXMPLR, QB=>OPEN, D
      =>nx25663, CLK=>clk, R=>rst);
   max_calc_reg_answer_11 : dffr port map ( Q=>answer_11_EXMPLR, QB=>OPEN, D
      =>nx25673, CLK=>clk, R=>rst);
   max_calc_reg_answer_12 : dffr port map ( Q=>answer_12_EXMPLR, QB=>OPEN, D
      =>nx25683, CLK=>clk, R=>rst);
   max_calc_reg_answer_13 : dffr port map ( Q=>answer_13_EXMPLR, QB=>OPEN, D
      =>nx25693, CLK=>clk, R=>rst);
   max_calc_reg_answer_14 : dffr port map ( Q=>answer_14_EXMPLR, QB=>OPEN, D
      =>nx25703, CLK=>clk, R=>rst);
   max_calc_reg_answer_15 : dffr port map ( Q=>answer_15_EXMPLR, QB=>OPEN, D
      =>nx25713, CLK=>clk, R=>rst);
   tri_mdr_data_out_176 : tri01 port map ( Y=>mdr_data_out(176), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_177 : tri01 port map ( Y=>mdr_data_out(177), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_178 : tri01 port map ( Y=>mdr_data_out(178), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_179 : tri01 port map ( Y=>mdr_data_out(179), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_180 : tri01 port map ( Y=>mdr_data_out(180), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_181 : tri01 port map ( Y=>mdr_data_out(181), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_182 : tri01 port map ( Y=>mdr_data_out(182), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_183 : tri01 port map ( Y=>mdr_data_out(183), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_184 : tri01 port map ( Y=>mdr_data_out(184), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_185 : tri01 port map ( Y=>mdr_data_out(185), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_186 : tri01 port map ( Y=>mdr_data_out(186), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_187 : tri01 port map ( Y=>mdr_data_out(187), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_188 : tri01 port map ( Y=>mdr_data_out(188), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_189 : tri01 port map ( Y=>mdr_data_out(189), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_190 : tri01 port map ( Y=>mdr_data_out(190), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_191 : tri01 port map ( Y=>mdr_data_out(191), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_192 : tri01 port map ( Y=>mdr_data_out(192), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_193 : tri01 port map ( Y=>mdr_data_out(193), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_194 : tri01 port map ( Y=>mdr_data_out(194), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_195 : tri01 port map ( Y=>mdr_data_out(195), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_196 : tri01 port map ( Y=>mdr_data_out(196), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_197 : tri01 port map ( Y=>mdr_data_out(197), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_198 : tri01 port map ( Y=>mdr_data_out(198), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_199 : tri01 port map ( Y=>mdr_data_out(199), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_200 : tri01 port map ( Y=>mdr_data_out(200), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_201 : tri01 port map ( Y=>mdr_data_out(201), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_202 : tri01 port map ( Y=>mdr_data_out(202), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_203 : tri01 port map ( Y=>mdr_data_out(203), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_204 : tri01 port map ( Y=>mdr_data_out(204), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_205 : tri01 port map ( Y=>mdr_data_out(205), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_206 : tri01 port map ( Y=>mdr_data_out(206), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_207 : tri01 port map ( Y=>mdr_data_out(207), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_208 : tri01 port map ( Y=>mdr_data_out(208), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_209 : tri01 port map ( Y=>mdr_data_out(209), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_210 : tri01 port map ( Y=>mdr_data_out(210), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_211 : tri01 port map ( Y=>mdr_data_out(211), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_212 : tri01 port map ( Y=>mdr_data_out(212), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_213 : tri01 port map ( Y=>mdr_data_out(213), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_214 : tri01 port map ( Y=>mdr_data_out(214), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_215 : tri01 port map ( Y=>mdr_data_out(215), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_216 : tri01 port map ( Y=>mdr_data_out(216), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_217 : tri01 port map ( Y=>mdr_data_out(217), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_218 : tri01 port map ( Y=>mdr_data_out(218), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_219 : tri01 port map ( Y=>mdr_data_out(219), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_220 : tri01 port map ( Y=>mdr_data_out(220), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_221 : tri01 port map ( Y=>mdr_data_out(221), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_222 : tri01 port map ( Y=>mdr_data_out(222), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_223 : tri01 port map ( Y=>mdr_data_out(223), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_224 : tri01 port map ( Y=>mdr_data_out(224), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_225 : tri01 port map ( Y=>mdr_data_out(225), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_226 : tri01 port map ( Y=>mdr_data_out(226), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_227 : tri01 port map ( Y=>mdr_data_out(227), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_228 : tri01 port map ( Y=>mdr_data_out(228), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_229 : tri01 port map ( Y=>mdr_data_out(229), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_230 : tri01 port map ( Y=>mdr_data_out(230), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_231 : tri01 port map ( Y=>mdr_data_out(231), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_232 : tri01 port map ( Y=>mdr_data_out(232), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_233 : tri01 port map ( Y=>mdr_data_out(233), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_234 : tri01 port map ( Y=>mdr_data_out(234), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_235 : tri01 port map ( Y=>mdr_data_out(235), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_236 : tri01 port map ( Y=>mdr_data_out(236), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_237 : tri01 port map ( Y=>mdr_data_out(237), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_238 : tri01 port map ( Y=>mdr_data_out(238), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_239 : tri01 port map ( Y=>mdr_data_out(239), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_240 : tri01 port map ( Y=>mdr_data_out(240), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_241 : tri01 port map ( Y=>mdr_data_out(241), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_242 : tri01 port map ( Y=>mdr_data_out(242), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_243 : tri01 port map ( Y=>mdr_data_out(243), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_244 : tri01 port map ( Y=>mdr_data_out(244), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_245 : tri01 port map ( Y=>mdr_data_out(245), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_246 : tri01 port map ( Y=>mdr_data_out(246), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_247 : tri01 port map ( Y=>mdr_data_out(247), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_248 : tri01 port map ( Y=>mdr_data_out(248), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_249 : tri01 port map ( Y=>mdr_data_out(249), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_250 : tri01 port map ( Y=>mdr_data_out(250), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_251 : tri01 port map ( Y=>mdr_data_out(251), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_252 : tri01 port map ( Y=>mdr_data_out(252), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_253 : tri01 port map ( Y=>mdr_data_out(253), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_254 : tri01 port map ( Y=>mdr_data_out(254), A=>nx25757, 
      E=>initiate);
   tri_mdr_data_out_255 : tri01 port map ( Y=>mdr_data_out(255), A=>nx25757, 
      E=>initiate);
   reg_enable_mdr_out : dffr port map ( Q=>enable_mdr_out, QB=>OPEN, D=>
      nx25753, CLK=>clk, R=>rst);
   ix25754 : mux21_ni port map ( Y=>nx25753, A0=>enable_mdr_out, A1=>nx190, 
      S0=>nx19296);
   ix19297 : nor03_2x port map ( Y=>nx19296, A0=>nx12895, A1=>nx56, A2=>
      nx34359);
   ix34360 : oai21 port map ( Y=>nx34359, A0=>nx25879, A1=>nx35101, B0=>
      nx868);
   reg_enable_mdr_in : dffr port map ( Q=>enable_mdr_in, QB=>OPEN, D=>
      nx25743, CLK=>clk, R=>rst);
   ix25744 : mux21_ni port map ( Y=>nx25743, A0=>nx19276, A1=>enable_mdr_in, 
      S0=>nx34365);
   ix34366 : nand03 port map ( Y=>nx34365, A0=>nx19266, A1=>nx26129, A2=>
      nx19236);
   ix19267 : oai21 port map ( Y=>nx19266, A0=>nx34399, A1=>nx34368, B0=>
      nx174);
   ix34369 : nor02ii port map ( Y=>nx34368, A0=>nx34403, A1=>sub_state(1));
   reg_enable_mar_in : dffr port map ( Q=>enable_mar_in, QB=>OPEN, D=>
      nx25733, CLK=>clk, R=>rst);
   ix25734 : mux21_ni port map ( Y=>nx25733, A0=>nx19250, A1=>enable_mar_in, 
      S0=>nx34377);
   ix19251 : ao22 port map ( Y=>nx19250, A0=>nx34403, A1=>nx174, B0=>nx12879, 
      B1=>nx26664);
   ix34378 : oai21 port map ( Y=>nx34377, A0=>nx35157, A1=>nx25916, B0=>
      nx19240);
   ix19233 : nor03_2x port map ( Y=>nx19232, A0=>nx258, A1=>nx12891, A2=>
      nx35155);
   ix19237 : inv01 port map ( Y=>nx19236, A=>nx34380);
   ix15325 : inv01 port map ( Y=>nx13370, A=>nx32050);
   ix15261 : inv01 port map ( Y=>nx13368, A=>nx32035);
   ix15197 : inv01 port map ( Y=>nx13365, A=>nx32020);
   ix15133 : inv01 port map ( Y=>nx13361, A=>nx32005);
   ix15069 : inv01 port map ( Y=>nx13359, A=>nx31990);
   ix15005 : inv01 port map ( Y=>nx13357, A=>nx31975);
   ix14941 : inv01 port map ( Y=>nx13355, A=>nx31961);
   ix31818 : inv01 port map ( Y=>nx31817, A=>nx14484);
   ix31811 : inv01 port map ( Y=>nx31810, A=>nx13351);
   ix14471 : inv01 port map ( Y=>nx14470, A=>nx31826);
   ix31816 : inv01 port map ( Y=>nx31815, A=>nx14460);
   ix14457 : inv01 port map ( Y=>nx14456, A=>nx31797);
   ix31783 : inv01 port map ( Y=>nx31782, A=>nx14436);
   ix31776 : inv01 port map ( Y=>nx31775, A=>nx13348);
   ix14423 : inv01 port map ( Y=>nx14422, A=>nx31829);
   ix31781 : inv01 port map ( Y=>nx31780, A=>nx14412);
   ix14409 : inv01 port map ( Y=>nx14408, A=>nx31762);
   ix31748 : inv01 port map ( Y=>nx31747, A=>nx14388);
   ix31741 : inv01 port map ( Y=>nx31740, A=>nx13346);
   ix14375 : inv01 port map ( Y=>nx14374, A=>nx31832);
   ix31746 : inv01 port map ( Y=>nx31745, A=>nx14364);
   ix14361 : inv01 port map ( Y=>nx14360, A=>nx31727);
   ix31713 : inv01 port map ( Y=>nx31712, A=>nx14340);
   ix31706 : inv01 port map ( Y=>nx31705, A=>nx13344);
   ix14327 : inv01 port map ( Y=>nx14326, A=>nx31835);
   ix31711 : inv01 port map ( Y=>nx31710, A=>nx14316);
   ix14313 : inv01 port map ( Y=>nx14312, A=>nx31692);
   ix31678 : inv01 port map ( Y=>nx31677, A=>nx14292);
   ix31671 : inv01 port map ( Y=>nx31670, A=>nx13341);
   ix14279 : inv01 port map ( Y=>nx14278, A=>nx31838);
   ix31676 : inv01 port map ( Y=>nx31675, A=>nx14268);
   ix14265 : inv01 port map ( Y=>nx14264, A=>nx31657);
   ix31643 : inv01 port map ( Y=>nx31642, A=>nx14244);
   ix31636 : inv01 port map ( Y=>nx31635, A=>nx13337);
   ix14231 : inv01 port map ( Y=>nx14230, A=>nx31841);
   ix31641 : inv01 port map ( Y=>nx31640, A=>nx14220);
   ix14217 : inv01 port map ( Y=>nx14216, A=>nx31618);
   ix31604 : inv01 port map ( Y=>nx31603, A=>nx14196);
   ix31599 : inv01 port map ( Y=>nx31598, A=>nx13335);
   ix14183 : inv01 port map ( Y=>nx14182, A=>nx31844);
   ix14009 : inv01 port map ( Y=>nx13332, A=>nx32239);
   ix13945 : inv01 port map ( Y=>nx13329, A=>nx32224);
   ix13881 : inv01 port map ( Y=>nx13325, A=>nx32209);
   ix13817 : inv01 port map ( Y=>nx13323, A=>nx32194);
   ix13753 : inv01 port map ( Y=>nx13321, A=>nx32179);
   ix13689 : inv01 port map ( Y=>nx13319, A=>nx32164);
   ix13625 : inv01 port map ( Y=>nx13315, A=>nx32150);
   ix31379 : inv01 port map ( Y=>nx31378, A=>nx13168);
   ix31372 : inv01 port map ( Y=>nx31371, A=>nx13312);
   ix13155 : inv01 port map ( Y=>nx13154, A=>nx31387);
   ix31377 : inv01 port map ( Y=>nx31376, A=>nx13144);
   ix13141 : inv01 port map ( Y=>nx13140, A=>nx31358);
   ix31344 : inv01 port map ( Y=>nx31343, A=>nx13120);
   ix31337 : inv01 port map ( Y=>nx31336, A=>nx13310);
   ix13107 : inv01 port map ( Y=>nx13106, A=>nx31390);
   ix31342 : inv01 port map ( Y=>nx31341, A=>nx13096);
   ix13093 : inv01 port map ( Y=>nx13092, A=>nx31323);
   ix31309 : inv01 port map ( Y=>nx31308, A=>nx13072);
   ix31302 : inv01 port map ( Y=>nx31301, A=>nx13308);
   ix13059 : inv01 port map ( Y=>nx13058, A=>nx31393);
   ix31307 : inv01 port map ( Y=>nx31306, A=>nx13048);
   ix13045 : inv01 port map ( Y=>nx13044, A=>nx31288);
   ix31274 : inv01 port map ( Y=>nx31273, A=>nx13024);
   ix31267 : inv01 port map ( Y=>nx31266, A=>nx13305);
   ix13011 : inv01 port map ( Y=>nx13010, A=>nx31396);
   ix31272 : inv01 port map ( Y=>nx31271, A=>nx13000);
   ix12997 : inv01 port map ( Y=>nx12996, A=>nx31253);
   ix31239 : inv01 port map ( Y=>nx31238, A=>nx12976);
   ix31232 : inv01 port map ( Y=>nx31231, A=>nx13301);
   ix12963 : inv01 port map ( Y=>nx12962, A=>nx31399);
   ix31237 : inv01 port map ( Y=>nx31236, A=>nx12952);
   ix12949 : inv01 port map ( Y=>nx12948, A=>nx31218);
   ix31204 : inv01 port map ( Y=>nx31203, A=>nx12928);
   ix31197 : inv01 port map ( Y=>nx31196, A=>nx13299);
   ix12915 : inv01 port map ( Y=>nx12914, A=>nx31402);
   ix31202 : inv01 port map ( Y=>nx31201, A=>nx12904);
   ix12901 : inv01 port map ( Y=>nx12900, A=>nx31179);
   ix31165 : inv01 port map ( Y=>nx31164, A=>nx12880);
   ix31160 : inv01 port map ( Y=>nx31159, A=>nx13297);
   ix12867 : inv01 port map ( Y=>nx12866, A=>nx31405);
   ix12141 : inv01 port map ( Y=>nx13293, A=>nx30123);
   ix12077 : inv01 port map ( Y=>nx13289, A=>nx30108);
   ix12013 : inv01 port map ( Y=>nx13287, A=>nx30093);
   ix11949 : inv01 port map ( Y=>nx13285, A=>nx30078);
   ix11885 : inv01 port map ( Y=>nx13283, A=>nx30063);
   ix11821 : inv01 port map ( Y=>nx13279, A=>nx30048);
   ix11757 : inv01 port map ( Y=>nx13276, A=>nx30034);
   ix29891 : inv01 port map ( Y=>nx29890, A=>nx11300);
   ix29884 : inv01 port map ( Y=>nx29883, A=>nx13274);
   ix11287 : inv01 port map ( Y=>nx11286, A=>nx29899);
   ix29889 : inv01 port map ( Y=>nx29888, A=>nx11276);
   ix11273 : inv01 port map ( Y=>nx11272, A=>nx29870);
   ix29856 : inv01 port map ( Y=>nx29855, A=>nx11252);
   ix29849 : inv01 port map ( Y=>nx29848, A=>nx13272);
   ix11239 : inv01 port map ( Y=>nx11238, A=>nx29902);
   ix29854 : inv01 port map ( Y=>nx29853, A=>nx11228);
   ix11225 : inv01 port map ( Y=>nx11224, A=>nx29835);
   ix29821 : inv01 port map ( Y=>nx29820, A=>nx11204);
   ix29814 : inv01 port map ( Y=>nx29813, A=>nx13269);
   ix11191 : inv01 port map ( Y=>nx11190, A=>nx29905);
   ix29819 : inv01 port map ( Y=>nx29818, A=>nx11180);
   ix11177 : inv01 port map ( Y=>nx11176, A=>nx29800);
   ix29786 : inv01 port map ( Y=>nx29785, A=>nx11156);
   ix29779 : inv01 port map ( Y=>nx29778, A=>nx13265);
   ix11143 : inv01 port map ( Y=>nx11142, A=>nx29908);
   ix29784 : inv01 port map ( Y=>nx29783, A=>nx11132);
   ix11129 : inv01 port map ( Y=>nx11128, A=>nx29765);
   ix29751 : inv01 port map ( Y=>nx29750, A=>nx11108);
   ix29744 : inv01 port map ( Y=>nx29743, A=>nx13263);
   ix11095 : inv01 port map ( Y=>nx11094, A=>nx29911);
   ix29749 : inv01 port map ( Y=>nx29748, A=>nx11084);
   ix11081 : inv01 port map ( Y=>nx11080, A=>nx29730);
   ix29716 : inv01 port map ( Y=>nx29715, A=>nx11060);
   ix29709 : inv01 port map ( Y=>nx29708, A=>nx13261);
   ix11047 : inv01 port map ( Y=>nx11046, A=>nx29914);
   ix29714 : inv01 port map ( Y=>nx29713, A=>nx11036);
   ix11033 : inv01 port map ( Y=>nx11032, A=>nx29691);
   ix29677 : inv01 port map ( Y=>nx29676, A=>nx11012);
   ix29672 : inv01 port map ( Y=>nx29671, A=>nx13259);
   ix10999 : inv01 port map ( Y=>nx10998, A=>nx29917);
   ix10819 : inv01 port map ( Y=>nx13253, A=>nx30312);
   ix10755 : inv01 port map ( Y=>nx13251, A=>nx30297);
   ix10691 : inv01 port map ( Y=>nx13249, A=>nx30282);
   ix10627 : inv01 port map ( Y=>nx13247, A=>nx30267);
   ix10563 : inv01 port map ( Y=>nx13243, A=>nx30252);
   ix10499 : inv01 port map ( Y=>nx13240, A=>nx30237);
   ix10435 : inv01 port map ( Y=>nx13238, A=>nx30223);
   ix29450 : inv01 port map ( Y=>nx29449, A=>nx9978);
   ix29443 : inv01 port map ( Y=>nx29442, A=>nx13236);
   ix9965 : inv01 port map ( Y=>nx9964, A=>nx29458);
   ix29448 : inv01 port map ( Y=>nx29447, A=>nx9954);
   ix9951 : inv01 port map ( Y=>nx9950, A=>nx29429);
   ix29415 : inv01 port map ( Y=>nx29414, A=>nx9930);
   ix29408 : inv01 port map ( Y=>nx29407, A=>nx13233);
   ix9917 : inv01 port map ( Y=>nx9916, A=>nx29461);
   ix29413 : inv01 port map ( Y=>nx29412, A=>nx9906);
   ix9903 : inv01 port map ( Y=>nx9902, A=>nx29394);
   ix29380 : inv01 port map ( Y=>nx29379, A=>nx9882);
   ix29373 : inv01 port map ( Y=>nx29372, A=>nx13229);
   ix9869 : inv01 port map ( Y=>nx9868, A=>nx29464);
   ix29378 : inv01 port map ( Y=>nx29377, A=>nx9858);
   ix9855 : inv01 port map ( Y=>nx9854, A=>nx29359);
   ix29345 : inv01 port map ( Y=>nx29344, A=>nx9834);
   ix29338 : inv01 port map ( Y=>nx29337, A=>nx13227);
   ix9821 : inv01 port map ( Y=>nx9820, A=>nx29467);
   ix29343 : inv01 port map ( Y=>nx29342, A=>nx9810);
   ix9807 : inv01 port map ( Y=>nx9806, A=>nx29324);
   ix29310 : inv01 port map ( Y=>nx29309, A=>nx9786);
   ix29303 : inv01 port map ( Y=>nx29302, A=>nx13225);
   ix9773 : inv01 port map ( Y=>nx9772, A=>nx29470);
   ix29308 : inv01 port map ( Y=>nx29307, A=>nx9762);
   ix9759 : inv01 port map ( Y=>nx9758, A=>nx29289);
   ix29275 : inv01 port map ( Y=>nx29274, A=>nx9738);
   ix29268 : inv01 port map ( Y=>nx29267, A=>nx13223);
   ix9725 : inv01 port map ( Y=>nx9724, A=>nx29473);
   ix29273 : inv01 port map ( Y=>nx29272, A=>nx9714);
   ix9711 : inv01 port map ( Y=>nx9710, A=>nx29250);
   ix29236 : inv01 port map ( Y=>nx29235, A=>nx9690);
   ix29231 : inv01 port map ( Y=>nx29230, A=>nx13219);
   ix9677 : inv01 port map ( Y=>nx9676, A=>nx29476);
   ix9011 : inv01 port map ( Y=>nx13215, A=>nx27943);
   ix8947 : inv01 port map ( Y=>nx13213, A=>nx27928);
   ix8883 : inv01 port map ( Y=>nx13211, A=>nx27913);
   ix8819 : inv01 port map ( Y=>nx13207, A=>nx27898);
   ix8755 : inv01 port map ( Y=>nx13204, A=>nx27883);
   ix8691 : inv01 port map ( Y=>nx13202, A=>nx27868);
   ix8627 : inv01 port map ( Y=>nx13200, A=>nx27854);
   ix8561 : inv01 port map ( Y=>nx13199, A=>nx27754);
   ix8497 : inv01 port map ( Y=>nx13195, A=>nx27739);
   ix8433 : inv01 port map ( Y=>nx13191, A=>nx27724);
   ix8369 : inv01 port map ( Y=>nx13187, A=>nx27709);
   ix8305 : inv01 port map ( Y=>nx13183, A=>nx27694);
   ix8241 : inv01 port map ( Y=>nx13179, A=>nx27679);
   ix8177 : inv01 port map ( Y=>nx13175, A=>nx27665);
   ix27522 : inv01 port map ( Y=>nx27521, A=>nx7720);
   ix27515 : inv01 port map ( Y=>nx27514, A=>nx13171);
   ix7707 : inv01 port map ( Y=>nx7706, A=>nx27530);
   ix27520 : inv01 port map ( Y=>nx27519, A=>nx7696);
   ix7693 : inv01 port map ( Y=>nx7692, A=>nx27501);
   ix27487 : inv01 port map ( Y=>nx27486, A=>nx7672);
   ix27480 : inv01 port map ( Y=>nx27479, A=>nx13169);
   ix7659 : inv01 port map ( Y=>nx7658, A=>nx27533);
   ix27485 : inv01 port map ( Y=>nx27484, A=>nx7648);
   ix7645 : inv01 port map ( Y=>nx7644, A=>nx27466);
   ix27452 : inv01 port map ( Y=>nx27451, A=>nx7624);
   ix27445 : inv01 port map ( Y=>nx27444, A=>nx13165);
   ix7611 : inv01 port map ( Y=>nx7610, A=>nx27536);
   ix27450 : inv01 port map ( Y=>nx27449, A=>nx7600);
   ix7597 : inv01 port map ( Y=>nx7596, A=>nx27431);
   ix27417 : inv01 port map ( Y=>nx27416, A=>nx7576);
   ix27410 : inv01 port map ( Y=>nx27409, A=>nx13162);
   ix7563 : inv01 port map ( Y=>nx7562, A=>nx27539);
   ix27415 : inv01 port map ( Y=>nx27414, A=>nx7552);
   ix7549 : inv01 port map ( Y=>nx7548, A=>nx27396);
   ix27382 : inv01 port map ( Y=>nx27381, A=>nx7528);
   ix27375 : inv01 port map ( Y=>nx27374, A=>nx13159);
   ix7515 : inv01 port map ( Y=>nx7514, A=>nx27542);
   ix27380 : inv01 port map ( Y=>nx27379, A=>nx7504);
   ix7501 : inv01 port map ( Y=>nx7500, A=>nx27361);
   ix27347 : inv01 port map ( Y=>nx27346, A=>nx7480);
   ix27340 : inv01 port map ( Y=>nx27339, A=>nx13155);
   ix7467 : inv01 port map ( Y=>nx7466, A=>nx27545);
   ix27345 : inv01 port map ( Y=>nx27344, A=>nx7456);
   ix7453 : inv01 port map ( Y=>nx7452, A=>nx27322);
   ix27308 : inv01 port map ( Y=>nx27307, A=>nx7432);
   ix27303 : inv01 port map ( Y=>nx27302, A=>nx13151);
   ix7419 : inv01 port map ( Y=>nx7418, A=>nx27548);
   ix27083 : inv01 port map ( Y=>nx27082, A=>nx6840);
   ix27076 : inv01 port map ( Y=>nx27075, A=>nx13146);
   ix6827 : inv01 port map ( Y=>nx6826, A=>nx27091);
   ix27081 : inv01 port map ( Y=>nx27080, A=>nx6816);
   ix6813 : inv01 port map ( Y=>nx6812, A=>nx27062);
   ix27048 : inv01 port map ( Y=>nx27047, A=>nx6792);
   ix27041 : inv01 port map ( Y=>nx27040, A=>nx13143);
   ix6779 : inv01 port map ( Y=>nx6778, A=>nx27094);
   ix27046 : inv01 port map ( Y=>nx27045, A=>nx6768);
   ix6765 : inv01 port map ( Y=>nx6764, A=>nx27027);
   ix27013 : inv01 port map ( Y=>nx27012, A=>nx6744);
   ix27006 : inv01 port map ( Y=>nx27005, A=>nx13139);
   ix6731 : inv01 port map ( Y=>nx6730, A=>nx27097);
   ix27011 : inv01 port map ( Y=>nx27010, A=>nx6720);
   ix6717 : inv01 port map ( Y=>nx6716, A=>nx26992);
   ix26978 : inv01 port map ( Y=>nx26977, A=>nx6696);
   ix26971 : inv01 port map ( Y=>nx26970, A=>nx13137);
   ix6683 : inv01 port map ( Y=>nx6682, A=>nx27100);
   ix26976 : inv01 port map ( Y=>nx26975, A=>nx6672);
   ix6669 : inv01 port map ( Y=>nx6668, A=>nx26957);
   ix26943 : inv01 port map ( Y=>nx26942, A=>nx6648);
   ix26936 : inv01 port map ( Y=>nx26935, A=>nx13133);
   ix6635 : inv01 port map ( Y=>nx6634, A=>nx27103);
   ix26941 : inv01 port map ( Y=>nx26940, A=>nx6624);
   ix6621 : inv01 port map ( Y=>nx6620, A=>nx26922);
   ix26908 : inv01 port map ( Y=>nx26907, A=>nx6600);
   ix26901 : inv01 port map ( Y=>nx26900, A=>nx13129);
   ix6587 : inv01 port map ( Y=>nx6586, A=>nx27106);
   ix26906 : inv01 port map ( Y=>nx26905, A=>nx6576);
   ix6573 : inv01 port map ( Y=>nx6572, A=>nx26883);
   ix26869 : inv01 port map ( Y=>nx26868, A=>nx6552);
   ix26864 : inv01 port map ( Y=>nx26863, A=>nx13125);
   ix6539 : inv01 port map ( Y=>nx6538, A=>nx27109);
   ix6353 : inv01 port map ( Y=>nx6352, A=>nx28172);
   ix6245 : inv01 port map ( Y=>nx6244, A=>nx26182);
   ix6181 : inv01 port map ( Y=>nx13114, A=>nx33671);
   ix6117 : inv01 port map ( Y=>nx13111, A=>nx33656);
   ix6053 : inv01 port map ( Y=>nx13107, A=>nx33641);
   ix5989 : inv01 port map ( Y=>nx13103, A=>nx33626);
   ix5925 : inv01 port map ( Y=>nx13099, A=>nx33611);
   ix5861 : inv01 port map ( Y=>nx13097, A=>nx33596);
   ix5797 : inv01 port map ( Y=>nx13093, A=>nx33582);
   ix26604 : inv01 port map ( Y=>nx26603, A=>nx5340);
   ix26597 : inv01 port map ( Y=>nx26596, A=>nx13090);
   ix5327 : inv01 port map ( Y=>nx5326, A=>nx26612);
   ix26602 : inv01 port map ( Y=>nx26601, A=>nx5316);
   ix5313 : inv01 port map ( Y=>nx5312, A=>nx26583);
   ix26569 : inv01 port map ( Y=>nx26568, A=>nx5292);
   ix26562 : inv01 port map ( Y=>nx26561, A=>nx13087);
   ix5279 : inv01 port map ( Y=>nx5278, A=>nx26615);
   ix26567 : inv01 port map ( Y=>nx26566, A=>nx5268);
   ix5265 : inv01 port map ( Y=>nx5264, A=>nx26548);
   ix26534 : inv01 port map ( Y=>nx26533, A=>nx5244);
   ix26527 : inv01 port map ( Y=>nx26526, A=>nx13083);
   ix5231 : inv01 port map ( Y=>nx5230, A=>nx26618);
   ix26532 : inv01 port map ( Y=>nx26531, A=>nx5220);
   ix5217 : inv01 port map ( Y=>nx5216, A=>nx26513);
   ix26499 : inv01 port map ( Y=>nx26498, A=>nx5196);
   ix26492 : inv01 port map ( Y=>nx26491, A=>nx13079);
   ix5183 : inv01 port map ( Y=>nx5182, A=>nx26621);
   ix26497 : inv01 port map ( Y=>nx26496, A=>nx5172);
   ix5169 : inv01 port map ( Y=>nx5168, A=>nx26478);
   ix26464 : inv01 port map ( Y=>nx26463, A=>nx5148);
   ix26457 : inv01 port map ( Y=>nx26456, A=>nx13075);
   ix5135 : inv01 port map ( Y=>nx5134, A=>nx26624);
   ix26462 : inv01 port map ( Y=>nx26461, A=>nx5124);
   ix5121 : inv01 port map ( Y=>nx5120, A=>nx26443);
   ix26429 : inv01 port map ( Y=>nx26428, A=>nx5100);
   ix26422 : inv01 port map ( Y=>nx26421, A=>nx13073);
   ix5087 : inv01 port map ( Y=>nx5086, A=>nx26627);
   ix26427 : inv01 port map ( Y=>nx26426, A=>nx5076);
   ix5073 : inv01 port map ( Y=>nx5072, A=>nx26404);
   ix26390 : inv01 port map ( Y=>nx26389, A=>nx5052);
   ix26385 : inv01 port map ( Y=>nx26384, A=>nx13069);
   ix5039 : inv01 port map ( Y=>nx5038, A=>nx26630);
   ix4843 : inv01 port map ( Y=>nx13063, A=>nx33473);
   ix4779 : inv01 port map ( Y=>nx13059, A=>nx33458);
   ix4715 : inv01 port map ( Y=>nx13055, A=>nx33443);
   ix4651 : inv01 port map ( Y=>nx13051, A=>nx33428);
   ix4587 : inv01 port map ( Y=>nx13049, A=>nx33413);
   ix4523 : inv01 port map ( Y=>nx13045, A=>nx33398);
   ix4459 : inv01 port map ( Y=>nx13042, A=>nx33384);
   ix28564 : inv01 port map ( Y=>nx28563, A=>nx4002);
   ix28557 : inv01 port map ( Y=>nx28556, A=>nx13039);
   ix3989 : inv01 port map ( Y=>nx3988, A=>nx28572);
   ix28562 : inv01 port map ( Y=>nx28561, A=>nx3978);
   ix3975 : inv01 port map ( Y=>nx3974, A=>nx28543);
   ix28529 : inv01 port map ( Y=>nx28528, A=>nx3954);
   ix28522 : inv01 port map ( Y=>nx28521, A=>nx13035);
   ix3941 : inv01 port map ( Y=>nx3940, A=>nx28575);
   ix28527 : inv01 port map ( Y=>nx28526, A=>nx3930);
   ix3927 : inv01 port map ( Y=>nx3926, A=>nx28508);
   ix28494 : inv01 port map ( Y=>nx28493, A=>nx3906);
   ix28487 : inv01 port map ( Y=>nx28486, A=>nx13031);
   ix3893 : inv01 port map ( Y=>nx3892, A=>nx28578);
   ix28492 : inv01 port map ( Y=>nx28491, A=>nx3882);
   ix3879 : inv01 port map ( Y=>nx3878, A=>nx28473);
   ix28459 : inv01 port map ( Y=>nx28458, A=>nx3858);
   ix28452 : inv01 port map ( Y=>nx28451, A=>nx13027);
   ix3845 : inv01 port map ( Y=>nx3844, A=>nx28581);
   ix28457 : inv01 port map ( Y=>nx28456, A=>nx3834);
   ix3831 : inv01 port map ( Y=>nx3830, A=>nx28438);
   ix28424 : inv01 port map ( Y=>nx28423, A=>nx3810);
   ix28417 : inv01 port map ( Y=>nx28416, A=>nx13025);
   ix3797 : inv01 port map ( Y=>nx3796, A=>nx28584);
   ix28422 : inv01 port map ( Y=>nx28421, A=>nx3786);
   ix3783 : inv01 port map ( Y=>nx3782, A=>nx28403);
   ix28389 : inv01 port map ( Y=>nx28388, A=>nx3762);
   ix28382 : inv01 port map ( Y=>nx28381, A=>nx13021);
   ix3749 : inv01 port map ( Y=>nx3748, A=>nx28587);
   ix28387 : inv01 port map ( Y=>nx28386, A=>nx3738);
   ix3735 : inv01 port map ( Y=>nx3734, A=>nx28364);
   ix28350 : inv01 port map ( Y=>nx28349, A=>nx3714);
   ix28345 : inv01 port map ( Y=>nx28344, A=>nx13018);
   ix3701 : inv01 port map ( Y=>nx3700, A=>nx28590);
   ix3505 : inv01 port map ( Y=>nx13011, A=>nx32850);
   ix3441 : inv01 port map ( Y=>nx13007, A=>nx32835);
   ix3377 : inv01 port map ( Y=>nx13003, A=>nx32820);
   ix3313 : inv01 port map ( Y=>nx13001, A=>nx32805);
   ix3249 : inv01 port map ( Y=>nx12997, A=>nx32790);
   ix3185 : inv01 port map ( Y=>nx12994, A=>nx32775);
   ix3121 : inv01 port map ( Y=>nx12991, A=>nx32761);
   ix29007 : inv01 port map ( Y=>nx29006, A=>nx2664);
   ix29000 : inv01 port map ( Y=>nx28999, A=>nx12987);
   ix2651 : inv01 port map ( Y=>nx2650, A=>nx29015);
   ix29005 : inv01 port map ( Y=>nx29004, A=>nx2640);
   ix2637 : inv01 port map ( Y=>nx2636, A=>nx28986);
   ix28972 : inv01 port map ( Y=>nx28971, A=>nx2616);
   ix28965 : inv01 port map ( Y=>nx28964, A=>nx12983);
   ix2603 : inv01 port map ( Y=>nx2602, A=>nx29018);
   ix28970 : inv01 port map ( Y=>nx28969, A=>nx2592);
   ix2589 : inv01 port map ( Y=>nx2588, A=>nx28951);
   ix28937 : inv01 port map ( Y=>nx28936, A=>nx2568);
   ix28930 : inv01 port map ( Y=>nx28929, A=>nx12979);
   ix2555 : inv01 port map ( Y=>nx2554, A=>nx29021);
   ix28935 : inv01 port map ( Y=>nx28934, A=>nx2544);
   ix2541 : inv01 port map ( Y=>nx2540, A=>nx28916);
   ix28902 : inv01 port map ( Y=>nx28901, A=>nx2520);
   ix28895 : inv01 port map ( Y=>nx28894, A=>nx12977);
   ix2507 : inv01 port map ( Y=>nx2506, A=>nx29024);
   ix28900 : inv01 port map ( Y=>nx28899, A=>nx2496);
   ix2493 : inv01 port map ( Y=>nx2492, A=>nx28881);
   ix28867 : inv01 port map ( Y=>nx28866, A=>nx2472);
   ix28860 : inv01 port map ( Y=>nx28859, A=>nx12973);
   ix2459 : inv01 port map ( Y=>nx2458, A=>nx29027);
   ix28865 : inv01 port map ( Y=>nx28864, A=>nx2448);
   ix2445 : inv01 port map ( Y=>nx2444, A=>nx28846);
   ix28832 : inv01 port map ( Y=>nx28831, A=>nx2424);
   ix28825 : inv01 port map ( Y=>nx28824, A=>nx12970);
   ix2411 : inv01 port map ( Y=>nx2410, A=>nx29030);
   ix28830 : inv01 port map ( Y=>nx28829, A=>nx2400);
   ix2397 : inv01 port map ( Y=>nx2396, A=>nx28807);
   ix28793 : inv01 port map ( Y=>nx28792, A=>nx2376);
   ix28788 : inv01 port map ( Y=>nx28787, A=>nx12967);
   ix2363 : inv01 port map ( Y=>nx2362, A=>nx29033);
   ix2167 : inv01 port map ( Y=>nx12959, A=>nx32654);
   ix2103 : inv01 port map ( Y=>nx12955, A=>nx32639);
   ix2039 : inv01 port map ( Y=>nx12953, A=>nx32624);
   ix1975 : inv01 port map ( Y=>nx12949, A=>nx32609);
   ix1911 : inv01 port map ( Y=>nx12946, A=>nx32594);
   ix1847 : inv01 port map ( Y=>nx12943, A=>nx32579);
   ix1783 : inv01 port map ( Y=>nx12939, A=>nx32565);
   ix30936 : inv01 port map ( Y=>nx30935, A=>nx1326);
   ix30929 : inv01 port map ( Y=>nx30928, A=>nx12935);
   ix1313 : inv01 port map ( Y=>nx1312, A=>nx30944);
   ix30934 : inv01 port map ( Y=>nx30933, A=>nx1302);
   ix1299 : inv01 port map ( Y=>nx1298, A=>nx30915);
   ix30901 : inv01 port map ( Y=>nx30900, A=>nx1278);
   ix30894 : inv01 port map ( Y=>nx30893, A=>nx12931);
   ix1265 : inv01 port map ( Y=>nx1264, A=>nx30947);
   ix30899 : inv01 port map ( Y=>nx30898, A=>nx1254);
   ix1251 : inv01 port map ( Y=>nx1250, A=>nx30880);
   ix30866 : inv01 port map ( Y=>nx30865, A=>nx1230);
   ix30859 : inv01 port map ( Y=>nx30858, A=>nx12929);
   ix1217 : inv01 port map ( Y=>nx1216, A=>nx30950);
   ix30864 : inv01 port map ( Y=>nx30863, A=>nx1206);
   ix1203 : inv01 port map ( Y=>nx1202, A=>nx30845);
   ix30831 : inv01 port map ( Y=>nx30830, A=>nx1182);
   ix30824 : inv01 port map ( Y=>nx30823, A=>nx12925);
   ix1169 : inv01 port map ( Y=>nx1168, A=>nx30953);
   ix30829 : inv01 port map ( Y=>nx30828, A=>nx1158);
   ix1155 : inv01 port map ( Y=>nx1154, A=>nx30810);
   ix30796 : inv01 port map ( Y=>nx30795, A=>nx1134);
   ix30789 : inv01 port map ( Y=>nx30788, A=>nx12922);
   ix1121 : inv01 port map ( Y=>nx1120, A=>nx30956);
   ix30794 : inv01 port map ( Y=>nx30793, A=>nx1110);
   ix1107 : inv01 port map ( Y=>nx1106, A=>nx30775);
   ix30761 : inv01 port map ( Y=>nx30760, A=>nx1086);
   ix30754 : inv01 port map ( Y=>nx30753, A=>nx12919);
   ix1073 : inv01 port map ( Y=>nx1072, A=>nx30959);
   ix30759 : inv01 port map ( Y=>nx30758, A=>nx1062);
   ix1059 : inv01 port map ( Y=>nx1058, A=>nx30736);
   ix30722 : inv01 port map ( Y=>nx30721, A=>nx1038);
   ix30717 : inv01 port map ( Y=>nx30716, A=>nx12915);
   ix1025 : inv01 port map ( Y=>nx1024, A=>nx30962);
   ix657 : inv01 port map ( Y=>nx656, A=>nx26056);
   ix549 : inv01 port map ( Y=>nx548, A=>nx26001);
   ix25836 : inv01 port map ( Y=>nx25835, A=>nx516);
   ix457 : inv01 port map ( Y=>nx12898, A=>nx25962);
   ix25920 : inv01 port map ( Y=>nx25919, A=>nx334);
   ix853 : inv01 port map ( Y=>nx12895, A=>nx26129);
   ix187 : inv01 port map ( Y=>nx186, A=>nx25907);
   ix25917 : inv01 port map ( Y=>nx25916, A=>nx174);
   ix25814 : inv01 port map ( Y=>nx25813, A=>nx12891);
   ix26665 : inv01 port map ( Y=>nx26664, A=>nx38);
   ix49 : inv01 port map ( Y=>nx12885, A=>nx25944);
   ix25901 : inv01 port map ( Y=>nx25900, A=>nx12879);
   ix34388 : inv02 port map ( Y=>nx34389, A=>nx35783);
   ix34390 : inv02 port map ( Y=>nx34391, A=>nx35783);
   ix34392 : inv02 port map ( Y=>nx34393, A=>nx35779);
   ix34394 : inv02 port map ( Y=>nx34395, A=>nx35779);
   ix34396 : inv02 port map ( Y=>nx34397, A=>nx35791);
   ix34398 : inv02 port map ( Y=>nx34399, A=>nx35791);
   ix34400 : buf02 port map ( Y=>nx34401, A=>sub_state(0));
   ix34402 : buf02 port map ( Y=>nx34403, A=>sub_state(0));
   ix34404 : inv02 port map ( Y=>nx34405, A=>nx35153);
   ix34406 : inv02 port map ( Y=>nx34407, A=>nx35153);
   ix34408 : inv02 port map ( Y=>nx34409, A=>nx35919);
   ix34418 : inv02 port map ( Y=>nx34419, A=>nx35925);
   ix34428 : inv02 port map ( Y=>nx34429, A=>nx35925);
   ix34456 : inv02 port map ( Y=>nx34457, A=>ready_signal);
   ix34458 : inv02 port map ( Y=>nx34459, A=>nx35589);
   ix34460 : inv02 port map ( Y=>nx34461, A=>nx35589);
   ix34462 : inv02 port map ( Y=>nx34463, A=>nx35589);
   ix34464 : inv02 port map ( Y=>nx34465, A=>nx35589);
   ix34466 : inv02 port map ( Y=>nx34467, A=>nx35589);
   ix34468 : inv02 port map ( Y=>nx34469, A=>nx35591);
   ix34470 : inv02 port map ( Y=>nx34471, A=>nx35591);
   ix34472 : inv02 port map ( Y=>nx34473, A=>nx35591);
   ix34474 : inv02 port map ( Y=>nx34475, A=>nx35591);
   ix34476 : inv02 port map ( Y=>nx34477, A=>nx35591);
   ix34478 : inv02 port map ( Y=>nx34479, A=>nx35591);
   ix34480 : inv02 port map ( Y=>nx34481, A=>nx35591);
   ix34482 : inv02 port map ( Y=>nx34483, A=>nx35593);
   ix34484 : inv02 port map ( Y=>nx34485, A=>nx35593);
   ix34486 : inv02 port map ( Y=>nx34487, A=>nx35593);
   ix34488 : inv02 port map ( Y=>nx34489, A=>nx35593);
   ix34490 : inv02 port map ( Y=>nx34491, A=>nx35593);
   ix34492 : inv02 port map ( Y=>nx34493, A=>nx35593);
   ix34494 : inv02 port map ( Y=>nx34495, A=>nx35101);
   ix34498 : inv02 port map ( Y=>nx34499, A=>nx25999);
   ix34500 : inv02 port map ( Y=>nx34501, A=>nx35799);
   ix34502 : buf02 port map ( Y=>nx34503, A=>enable_address);
   ix34504 : buf02 port map ( Y=>nx34505, A=>enable_address);
   ix34506 : buf02 port map ( Y=>nx34507, A=>nx350);
   ix34508 : buf02 port map ( Y=>nx34509, A=>nx350);
   ix34510 : inv02 port map ( Y=>nx34511, A=>nx35263);
   ix34512 : inv02 port map ( Y=>nx34513, A=>nx35265);
   ix34514 : inv02 port map ( Y=>nx34515, A=>nx35265);
   ix34516 : inv02 port map ( Y=>nx34517, A=>nx35265);
   ix34518 : inv02 port map ( Y=>nx34519, A=>nx35265);
   ix34520 : inv02 port map ( Y=>nx34521, A=>nx35265);
   ix34522 : inv02 port map ( Y=>nx34523, A=>nx35265);
   ix34524 : inv02 port map ( Y=>nx34525, A=>nx35265);
   ix34526 : inv02 port map ( Y=>nx34527, A=>nx35267);
   ix34528 : inv02 port map ( Y=>nx34529, A=>nx35267);
   ix34530 : inv02 port map ( Y=>nx34531, A=>nx35267);
   ix34532 : inv02 port map ( Y=>nx34533, A=>nx35267);
   ix34534 : inv02 port map ( Y=>nx34535, A=>nx35267);
   ix34536 : inv02 port map ( Y=>nx34537, A=>nx35267);
   ix34538 : inv02 port map ( Y=>nx34539, A=>nx35267);
   ix34540 : inv02 port map ( Y=>nx34541, A=>nx35269);
   ix34542 : inv02 port map ( Y=>nx34543, A=>nx35269);
   ix34544 : inv02 port map ( Y=>nx34545, A=>nx35269);
   ix34546 : inv02 port map ( Y=>nx34547, A=>nx35269);
   ix34548 : inv02 port map ( Y=>nx34549, A=>nx35269);
   ix34550 : inv02 port map ( Y=>nx34551, A=>nx35269);
   ix34552 : inv02 port map ( Y=>nx34553, A=>nx35269);
   ix34554 : inv02 port map ( Y=>nx34555, A=>nx35271);
   ix34556 : inv02 port map ( Y=>nx34557, A=>nx36147);
   ix34570 : inv02 port map ( Y=>nx34571, A=>nx36155);
   ix34578 : inv02 port map ( Y=>nx34579, A=>nx30744);
   ix34580 : inv02 port map ( Y=>nx34581, A=>nx30744);
   ix34582 : inv02 port map ( Y=>nx34583, A=>nx30744);
   ix34588 : inv02 port map ( Y=>nx34589, A=>nx36093);
   ix34602 : inv02 port map ( Y=>nx34603, A=>nx36101);
   ix34610 : inv02 port map ( Y=>nx34611, A=>nx28815);
   ix34612 : inv02 port map ( Y=>nx34613, A=>nx28815);
   ix34614 : inv02 port map ( Y=>nx34615, A=>nx28815);
   ix34620 : inv02 port map ( Y=>nx34621, A=>nx36077);
   ix34634 : inv02 port map ( Y=>nx34635, A=>nx36085);
   ix34642 : inv02 port map ( Y=>nx34643, A=>nx28372);
   ix34644 : inv02 port map ( Y=>nx34645, A=>nx28372);
   ix34646 : inv02 port map ( Y=>nx34647, A=>nx28372);
   ix34652 : inv02 port map ( Y=>nx34653, A=>nx36003);
   ix34666 : inv02 port map ( Y=>nx34667, A=>nx36011);
   ix34674 : inv02 port map ( Y=>nx34675, A=>nx26412);
   ix34676 : inv02 port map ( Y=>nx34677, A=>nx26412);
   ix34678 : inv02 port map ( Y=>nx34679, A=>nx26412);
   ix34704 : inv02 port map ( Y=>nx34705, A=>nx35977);
   ix34736 : inv02 port map ( Y=>nx34737, A=>nx34735);
   ix34738 : inv02 port map ( Y=>nx34739, A=>nx35843);
   ix34740 : inv02 port map ( Y=>nx34741, A=>nx35843);
   ix34742 : inv02 port map ( Y=>nx34743, A=>nx35843);
   ix34744 : inv02 port map ( Y=>nx34745, A=>nx35843);
   ix34746 : inv02 port map ( Y=>nx34747, A=>nx35361);
   ix34748 : inv02 port map ( Y=>nx34749, A=>nx35361);
   ix34750 : inv02 port map ( Y=>nx34751, A=>nx35361);
   ix34752 : inv02 port map ( Y=>nx34753, A=>nx36063);
   ix34754 : inv02 port map ( Y=>nx34755, A=>nx36063);
   ix34756 : inv02 port map ( Y=>nx34757, A=>nx36063);
   ix34758 : inv02 port map ( Y=>nx34759, A=>nx36063);
   ix34760 : inv02 port map ( Y=>nx34761, A=>nx36063);
   ix34762 : inv02 port map ( Y=>nx34763, A=>nx36063);
   ix34764 : inv02 port map ( Y=>nx34765, A=>nx36063);
   ix34766 : inv02 port map ( Y=>nx34767, A=>nx36067);
   ix34768 : inv02 port map ( Y=>nx34769, A=>nx36067);
   ix34770 : inv02 port map ( Y=>nx34771, A=>nx36067);
   ix34772 : inv02 port map ( Y=>nx34773, A=>nx36067);
   ix34774 : inv02 port map ( Y=>nx34775, A=>nx36067);
   ix34776 : inv02 port map ( Y=>nx34777, A=>nx36067);
   ix34778 : inv02 port map ( Y=>nx34779, A=>nx36067);
   ix34780 : inv02 port map ( Y=>nx34781, A=>nx36071);
   ix34782 : inv02 port map ( Y=>nx34783, A=>nx36071);
   ix34784 : inv02 port map ( Y=>nx34785, A=>nx36071);
   ix34786 : inv02 port map ( Y=>nx34787, A=>nx36071);
   ix34788 : inv02 port map ( Y=>nx34789, A=>nx36071);
   ix34790 : inv02 port map ( Y=>nx34791, A=>nx36071);
   ix34792 : inv02 port map ( Y=>nx34793, A=>nx36071);
   ix34794 : inv02 port map ( Y=>nx34795, A=>nx36075);
   ix34796 : inv02 port map ( Y=>nx34797, A=>nx36075);
   ix34798 : inv02 port map ( Y=>nx34799, A=>nx36075);
   ix34800 : inv02 port map ( Y=>nx34801, A=>nx36075);
   ix34802 : inv02 port map ( Y=>nx34803, A=>nx36075);
   ix34804 : inv02 port map ( Y=>nx34805, A=>nx36075);
   ix34806 : inv02 port map ( Y=>nx34807, A=>nx36075);
   ix34808 : inv02 port map ( Y=>nx34809, A=>nx35371);
   ix34810 : inv02 port map ( Y=>nx34811, A=>nx35371);
   ix34812 : inv02 port map ( Y=>nx34813, A=>nx35371);
   ix34814 : inv02 port map ( Y=>nx34815, A=>nx35371);
   ix34816 : inv02 port map ( Y=>nx34817, A=>nx35371);
   ix34818 : inv02 port map ( Y=>nx34819, A=>nx35371);
   ix34832 : inv02 port map ( Y=>nx34833, A=>nx36031);
   ix34846 : inv02 port map ( Y=>nx34847, A=>nx36039);
   ix34854 : inv02 port map ( Y=>nx34855, A=>nx26891);
   ix34856 : inv02 port map ( Y=>nx34857, A=>nx26891);
   ix34858 : inv02 port map ( Y=>nx34859, A=>nx26891);
   ix34864 : inv02 port map ( Y=>nx34865, A=>nx36047);
   ix34878 : inv02 port map ( Y=>nx34879, A=>nx36055);
   ix34886 : inv02 port map ( Y=>nx34887, A=>nx27330);
   ix34888 : inv02 port map ( Y=>nx34889, A=>nx27330);
   ix34890 : inv02 port map ( Y=>nx34891, A=>nx27330);
   ix34924 : inv02 port map ( Y=>nx34925, A=>nx36109);
   ix34938 : inv02 port map ( Y=>nx34939, A=>nx36117);
   ix34946 : inv02 port map ( Y=>nx34947, A=>nx29258);
   ix34948 : inv02 port map ( Y=>nx34949, A=>nx29258);
   ix34950 : inv02 port map ( Y=>nx34951, A=>nx29258);
   ix34956 : inv02 port map ( Y=>nx34957, A=>nx36131);
   ix34970 : inv02 port map ( Y=>nx34971, A=>nx36139);
   ix34978 : inv02 port map ( Y=>nx34979, A=>nx29699);
   ix34980 : inv02 port map ( Y=>nx34981, A=>nx29699);
   ix34982 : inv02 port map ( Y=>nx34983, A=>nx29699);
   ix34996 : inv02 port map ( Y=>nx34997, A=>nx36163);
   ix35010 : inv02 port map ( Y=>nx35011, A=>nx36171);
   ix35018 : inv02 port map ( Y=>nx35019, A=>nx31187);
   ix35020 : inv02 port map ( Y=>nx35021, A=>nx31187);
   ix35022 : inv02 port map ( Y=>nx35023, A=>nx31187);
   ix35028 : inv02 port map ( Y=>nx35029, A=>nx36179);
   ix35042 : inv02 port map ( Y=>nx35043, A=>nx36187);
   ix35050 : inv02 port map ( Y=>nx35051, A=>nx31626);
   ix35052 : inv02 port map ( Y=>nx35053, A=>nx31626);
   ix35054 : inv02 port map ( Y=>nx35055, A=>nx31626);
   ix35094 : buf02 port map ( Y=>nx35095, A=>nx25827);
   ix35096 : buf02 port map ( Y=>nx35097, A=>nx25827);
   ix35098 : inv02 port map ( Y=>nx35099, A=>nx12893);
   ix35100 : inv02 port map ( Y=>nx35101, A=>nx12893);
   ix35102 : inv02 port map ( Y=>nx35103, A=>nx36201);
   ix35148 : inv02 port map ( Y=>nx35149, A=>nx4);
   ix35152 : inv02 port map ( Y=>nx35153, A=>nx35713);
   ix35154 : inv02 port map ( Y=>nx35155, A=>nx12882);
   ix35156 : buf02 port map ( Y=>nx35157, A=>nx25896);
   ix35158 : buf02 port map ( Y=>nx35159, A=>nx25937);
   ix35160 : buf02 port map ( Y=>nx35161, A=>nx25937);
   ix35162 : inv02 port map ( Y=>nx35163, A=>enable_decoder_dst_booth);
   ix35164 : inv02 port map ( Y=>nx35165, A=>nx36307);
   ix35166 : inv02 port map ( Y=>nx35167, A=>nx36307);
   ix35168 : inv02 port map ( Y=>nx35169, A=>nx36307);
   ix35170 : inv02 port map ( Y=>nx35171, A=>nx36307);
   ix35172 : inv02 port map ( Y=>nx35173, A=>max_calc_state_2);
   ix35174 : inv02 port map ( Y=>nx35175, A=>nx36299);
   ix35176 : inv02 port map ( Y=>nx35177, A=>nx36299);
   ix35178 : inv02 port map ( Y=>nx35179, A=>nx36299);
   ix35180 : inv02 port map ( Y=>nx35181, A=>nx36299);
   ix35182 : inv02 port map ( Y=>nx35183, A=>nx36299);
   ix35184 : inv02 port map ( Y=>nx35185, A=>nx36299);
   ix35186 : inv02 port map ( Y=>nx35187, A=>max_calc_state_1);
   ix35188 : inv02 port map ( Y=>nx35189, A=>nx36331);
   ix35190 : inv02 port map ( Y=>nx35191, A=>nx36331);
   ix35192 : inv02 port map ( Y=>nx35193, A=>
      booth_booth_integrtaion_0_shift_reg_output_9);
   ix35194 : inv02 port map ( Y=>nx35195, A=>nx36327);
   ix35196 : inv02 port map ( Y=>nx35197, A=>nx36327);
   ix35198 : inv02 port map ( Y=>nx35199, A=>nx36327);
   ix35200 : inv01 port map ( Y=>nx35201, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix35204 : buf02 port map ( Y=>nx35205, A=>nx26386);
   ix35206 : buf02 port map ( Y=>nx35207, A=>nx26423);
   ix35208 : buf02 port map ( Y=>nx35209, A=>nx26458);
   ix35210 : buf02 port map ( Y=>nx35211, A=>nx26493);
   ix35212 : buf02 port map ( Y=>nx35213, A=>nx26528);
   ix35214 : buf02 port map ( Y=>nx35215, A=>nx26563);
   ix35216 : buf02 port map ( Y=>nx35217, A=>nx26598);
   ix35262 : inv02 port map ( Y=>nx35263, A=>nx36277);
   ix35264 : inv02 port map ( Y=>nx35265, A=>nx36277);
   ix35266 : inv02 port map ( Y=>nx35267, A=>nx36277);
   ix35268 : inv02 port map ( Y=>nx35269, A=>nx36277);
   ix35270 : inv02 port map ( Y=>nx35271, A=>nx36277);
   ix35300 : inv02 port map ( Y=>nx35301, A=>
      booth_booth_integrtaion_8_shift_reg_output_9);
   ix35302 : inv02 port map ( Y=>nx35303, A=>nx36341);
   ix35304 : inv02 port map ( Y=>nx35305, A=>nx36341);
   ix35306 : inv02 port map ( Y=>nx35307, A=>nx36341);
   ix35308 : inv01 port map ( Y=>nx35309, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix35312 : buf02 port map ( Y=>nx35313, A=>nx26865);
   ix35314 : buf02 port map ( Y=>nx35315, A=>nx26902);
   ix35316 : buf02 port map ( Y=>nx35317, A=>nx26937);
   ix35318 : buf02 port map ( Y=>nx35319, A=>nx26972);
   ix35320 : buf02 port map ( Y=>nx35321, A=>nx27007);
   ix35322 : buf02 port map ( Y=>nx35323, A=>nx27042);
   ix35324 : buf02 port map ( Y=>nx35325, A=>nx27077);
   ix35326 : inv02 port map ( Y=>nx35327, A=>
      booth_booth_integrtaion_9_shift_reg_output_9);
   ix35328 : inv02 port map ( Y=>nx35329, A=>nx36345);
   ix35330 : inv02 port map ( Y=>nx35331, A=>nx36345);
   ix35332 : inv02 port map ( Y=>nx35333, A=>nx36345);
   ix35334 : inv01 port map ( Y=>nx35335, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix35338 : buf02 port map ( Y=>nx35339, A=>nx27304);
   ix35340 : buf02 port map ( Y=>nx35341, A=>nx27341);
   ix35342 : buf02 port map ( Y=>nx35343, A=>nx27376);
   ix35344 : buf02 port map ( Y=>nx35345, A=>nx27411);
   ix35346 : buf02 port map ( Y=>nx35347, A=>nx27446);
   ix35348 : buf02 port map ( Y=>nx35349, A=>nx27481);
   ix35350 : buf02 port map ( Y=>nx35351, A=>nx27516);
   ix35360 : inv02 port map ( Y=>nx35361, A=>nx36281);
   ix35362 : inv02 port map ( Y=>nx35363, A=>nx36337);
   ix35364 : inv02 port map ( Y=>nx35365, A=>nx36337);
   ix35366 : inv02 port map ( Y=>nx35367, A=>nx36337);
   ix35368 : inv02 port map ( Y=>nx35369, A=>nx36337);
   ix35370 : inv02 port map ( Y=>nx35371, A=>nx36337);
   ix35372 : inv02 port map ( Y=>nx35373, A=>
      booth_booth_integrtaion_1_shift_reg_output_9);
   ix35374 : inv02 port map ( Y=>nx35375, A=>nx36323);
   ix35376 : inv02 port map ( Y=>nx35377, A=>nx36323);
   ix35378 : inv02 port map ( Y=>nx35379, A=>nx36323);
   ix35380 : inv01 port map ( Y=>nx35381, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix35384 : buf02 port map ( Y=>nx35385, A=>nx28346);
   ix35386 : buf02 port map ( Y=>nx35387, A=>nx28383);
   ix35388 : buf02 port map ( Y=>nx35389, A=>nx28418);
   ix35390 : buf02 port map ( Y=>nx35391, A=>nx28453);
   ix35392 : buf02 port map ( Y=>nx35393, A=>nx28488);
   ix35394 : buf02 port map ( Y=>nx35395, A=>nx28523);
   ix35396 : buf02 port map ( Y=>nx35397, A=>nx28558);
   ix35398 : inv02 port map ( Y=>nx35399, A=>
      booth_booth_integrtaion_2_shift_reg_output_9);
   ix35400 : inv02 port map ( Y=>nx35401, A=>nx36319);
   ix35402 : inv02 port map ( Y=>nx35403, A=>nx36319);
   ix35404 : inv02 port map ( Y=>nx35405, A=>nx36319);
   ix35406 : inv01 port map ( Y=>nx35407, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix35410 : buf02 port map ( Y=>nx35411, A=>nx28789);
   ix35412 : buf02 port map ( Y=>nx35413, A=>nx28826);
   ix35414 : buf02 port map ( Y=>nx35415, A=>nx28861);
   ix35416 : buf02 port map ( Y=>nx35417, A=>nx28896);
   ix35418 : buf02 port map ( Y=>nx35419, A=>nx28931);
   ix35420 : buf02 port map ( Y=>nx35421, A=>nx28966);
   ix35422 : buf02 port map ( Y=>nx35423, A=>nx29001);
   ix35424 : inv02 port map ( Y=>nx35425, A=>
      booth_booth_integrtaion_4_shift_reg_output_9);
   ix35426 : inv02 port map ( Y=>nx35427, A=>nx36349);
   ix35428 : inv02 port map ( Y=>nx35429, A=>nx36349);
   ix35430 : inv02 port map ( Y=>nx35431, A=>nx36349);
   ix35432 : inv01 port map ( Y=>nx35433, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix35436 : buf02 port map ( Y=>nx35437, A=>nx29232);
   ix35438 : buf02 port map ( Y=>nx35439, A=>nx29269);
   ix35440 : buf02 port map ( Y=>nx35441, A=>nx29304);
   ix35442 : buf02 port map ( Y=>nx35443, A=>nx29339);
   ix35444 : buf02 port map ( Y=>nx35445, A=>nx29374);
   ix35446 : buf02 port map ( Y=>nx35447, A=>nx29409);
   ix35448 : buf02 port map ( Y=>nx35449, A=>nx29444);
   ix35452 : inv02 port map ( Y=>nx35453, A=>nx36195);
   ix35454 : inv02 port map ( Y=>nx35455, A=>nx36195);
   ix35456 : inv02 port map ( Y=>nx35457, A=>nx36195);
   ix35458 : inv02 port map ( Y=>nx35459, A=>nx36195);
   ix35460 : inv02 port map ( Y=>nx35461, A=>nx36195);
   ix35462 : inv02 port map ( Y=>nx35463, A=>nx36125);
   ix35464 : inv02 port map ( Y=>nx35465, A=>nx36125);
   ix35466 : inv02 port map ( Y=>nx35467, A=>nx36125);
   ix35468 : inv02 port map ( Y=>nx35469, A=>nx36125);
   ix35472 : inv02 port map ( Y=>nx35473, A=>
      booth_booth_integrtaion_5_shift_reg_output_9);
   ix35474 : inv02 port map ( Y=>nx35475, A=>nx36353);
   ix35476 : inv02 port map ( Y=>nx35477, A=>nx36353);
   ix35478 : inv02 port map ( Y=>nx35479, A=>nx36353);
   ix35480 : inv01 port map ( Y=>nx35481, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix35484 : buf02 port map ( Y=>nx35485, A=>nx29673);
   ix35486 : buf02 port map ( Y=>nx35487, A=>nx29710);
   ix35488 : buf02 port map ( Y=>nx35489, A=>nx29745);
   ix35490 : buf02 port map ( Y=>nx35491, A=>nx29780);
   ix35492 : buf02 port map ( Y=>nx35493, A=>nx29815);
   ix35494 : buf02 port map ( Y=>nx35495, A=>nx29850);
   ix35496 : buf02 port map ( Y=>nx35497, A=>nx29885);
   ix35498 : inv02 port map ( Y=>nx35499, A=>
      booth_booth_integrtaion_3_shift_reg_output_9);
   ix35500 : inv02 port map ( Y=>nx35501, A=>nx36315);
   ix35502 : inv02 port map ( Y=>nx35503, A=>nx36315);
   ix35504 : inv02 port map ( Y=>nx35505, A=>nx36315);
   ix35506 : inv01 port map ( Y=>nx35507, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix35510 : buf02 port map ( Y=>nx35511, A=>nx30718);
   ix35512 : buf02 port map ( Y=>nx35513, A=>nx30755);
   ix35514 : buf02 port map ( Y=>nx35515, A=>nx30790);
   ix35516 : buf02 port map ( Y=>nx35517, A=>nx30825);
   ix35518 : buf02 port map ( Y=>nx35519, A=>nx30860);
   ix35520 : buf02 port map ( Y=>nx35521, A=>nx30895);
   ix35522 : buf02 port map ( Y=>nx35523, A=>nx30930);
   ix35524 : inv02 port map ( Y=>nx35525, A=>
      booth_booth_integrtaion_6_shift_reg_output_9);
   ix35526 : inv02 port map ( Y=>nx35527, A=>nx36357);
   ix35528 : inv02 port map ( Y=>nx35529, A=>nx36357);
   ix35530 : inv02 port map ( Y=>nx35531, A=>nx36357);
   ix35532 : inv01 port map ( Y=>nx35533, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix35536 : buf02 port map ( Y=>nx35537, A=>nx31161);
   ix35538 : buf02 port map ( Y=>nx35539, A=>nx31198);
   ix35540 : buf02 port map ( Y=>nx35541, A=>nx31233);
   ix35542 : buf02 port map ( Y=>nx35543, A=>nx31268);
   ix35544 : buf02 port map ( Y=>nx35545, A=>nx31303);
   ix35546 : buf02 port map ( Y=>nx35547, A=>nx31338);
   ix35548 : buf02 port map ( Y=>nx35549, A=>nx31373);
   ix35550 : inv02 port map ( Y=>nx35551, A=>
      booth_booth_integrtaion_7_shift_reg_output_9);
   ix35552 : inv02 port map ( Y=>nx35553, A=>nx36361);
   ix35554 : inv02 port map ( Y=>nx35555, A=>nx36361);
   ix35556 : inv02 port map ( Y=>nx35557, A=>nx36361);
   ix35558 : inv01 port map ( Y=>nx35559, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix35562 : buf02 port map ( Y=>nx35563, A=>nx31600);
   ix35564 : buf02 port map ( Y=>nx35565, A=>nx31637);
   ix35566 : buf02 port map ( Y=>nx35567, A=>nx31672);
   ix35568 : buf02 port map ( Y=>nx35569, A=>nx31707);
   ix35570 : buf02 port map ( Y=>nx35571, A=>nx31742);
   ix35572 : buf02 port map ( Y=>nx35573, A=>nx31777);
   ix35574 : buf02 port map ( Y=>nx35575, A=>nx31812);
   ix35588 : inv02 port map ( Y=>nx35589, A=>nx34457);
   ix35590 : inv02 port map ( Y=>nx35591, A=>nx34457);
   ix35592 : inv02 port map ( Y=>nx35593, A=>nx34457);
   ix35594 : inv02 port map ( Y=>nx35595, A=>nx25854);
   ix35596 : inv02 port map ( Y=>nx35597, A=>nx36365);
   ix35598 : inv02 port map ( Y=>nx35599, A=>nx36365);
   ix35600 : inv02 port map ( Y=>nx35601, A=>nx36365);
   ix35602 : inv02 port map ( Y=>nx35603, A=>nx26669);
   ix35604 : inv02 port map ( Y=>nx35605, A=>nx36373);
   ix35606 : inv02 port map ( Y=>nx35607, A=>nx36373);
   ix35608 : inv02 port map ( Y=>nx35609, A=>nx36373);
   ix35614 : inv02 port map ( Y=>nx35615, A=>ready_signal);
   ix13624 : nand02 port map ( Y=>nx13623, A0=>nx35911, A1=>nx35919);
   ix13614 : mux21_ni port map ( Y=>nx13613, A0=>nx34409, A1=>
      booth_shift_Reg_adder_0_output_17, S0=>nx35911);
   ix13604 : mux21_ni port map ( Y=>nx13603, A0=>
      booth_shift_Reg_adder_0_output_17, A1=>
      booth_shift_Reg_adder_0_output_16, S0=>nx35911);
   ix13594 : mux21_ni port map ( Y=>nx13593, A0=>
      booth_shift_Reg_adder_0_output_16, A1=>
      booth_shift_Reg_adder_0_output_15, S0=>nx35911);
   ix13584 : mux21_ni port map ( Y=>nx13583, A0=>
      booth_shift_Reg_adder_0_output_15, A1=>
      booth_shift_Reg_adder_0_output_14, S0=>nx35911);
   ix13574 : mux21_ni port map ( Y=>nx13573, A0=>
      booth_shift_Reg_adder_0_output_14, A1=>
      booth_shift_Reg_adder_0_output_13, S0=>nx35911);
   ix13564 : mux21_ni port map ( Y=>nx13563, A0=>
      booth_shift_Reg_adder_0_output_13, A1=>
      booth_shift_Reg_adder_0_output_12, S0=>nx35911);
   ix13554 : mux21_ni port map ( Y=>nx13553, A0=>
      booth_shift_Reg_adder_0_output_12, A1=>
      booth_shift_Reg_adder_0_output_11, S0=>nx35913);
   ix13544 : mux21_ni port map ( Y=>nx13543, A0=>
      booth_shift_Reg_adder_0_output_11, A1=>
      booth_shift_Reg_adder_0_output_10, S0=>nx35913);
   ix13534 : mux21_ni port map ( Y=>nx13533, A0=>
      booth_shift_Reg_adder_0_output_10, A1=>
      booth_shift_Reg_adder_0_output_9, S0=>nx35913);
   ix13524 : mux21_ni port map ( Y=>nx13523, A0=>
      booth_shift_Reg_adder_0_output_9, A1=>booth_shift_Reg_adder_0_output_8, 
      S0=>nx35913);
   ix13514 : mux21_ni port map ( Y=>nx13513, A0=>
      booth_shift_Reg_adder_0_output_8, A1=>booth_shift_Reg_adder_0_output_7, 
      S0=>nx35913);
   ix13504 : mux21_ni port map ( Y=>nx13503, A0=>
      booth_shift_Reg_adder_0_output_7, A1=>booth_shift_Reg_adder_0_output_6, 
      S0=>nx35913);
   ix13494 : mux21_ni port map ( Y=>nx13493, A0=>
      booth_shift_Reg_adder_0_output_6, A1=>booth_shift_Reg_adder_0_output_5, 
      S0=>nx35913);
   ix13484 : mux21_ni port map ( Y=>nx13483, A0=>
      booth_shift_Reg_adder_0_output_5, A1=>booth_shift_Reg_adder_0_output_4, 
      S0=>nx35915);
   ix13474 : mux21_ni port map ( Y=>nx13473, A0=>
      booth_shift_Reg_adder_0_output_4, A1=>booth_shift_Reg_adder_0_output_3, 
      S0=>nx35915);
   ix13464 : mux21_ni port map ( Y=>nx13463, A0=>
      booth_shift_Reg_adder_0_output_3, A1=>booth_shift_Reg_adder_0_output_2, 
      S0=>nx35915);
   ix13454 : mux21_ni port map ( Y=>nx13453, A0=>
      booth_shift_Reg_adder_0_output_2, A1=>booth_shift_Reg_adder_0_output_1, 
      S0=>nx35915);
   ix13444 : mux21_ni port map ( Y=>nx13443, A0=>
      booth_shift_Reg_adder_0_output_1, A1=>booth_shift_Reg_adder_0_output_0, 
      S0=>nx35915);
   ix13430 : nor02ii port map ( Y=>nx13429, A0=>nx35915, A1=>
      booth_shift_Reg_adder_0_output_0);
   ix13424 : mux21 port map ( Y=>nx13423, A0=>nx34457, A1=>nx35153, S0=>nx64
   );
   ix831 : ao221 port map ( Y=>nx830, A0=>nx35791, A1=>nx172, B0=>nx25944, 
      B1=>nx35713, C0=>nx35621);
   ix13634 : ao32 port map ( Y=>nx13633, A0=>nx35783, A1=>nx35779, A2=>
      nx25907, B0=>sub_state(2), B1=>nx35623);
   ix35622 : inv01 port map ( Y=>nx35623, A=>nx12883);
   ix14094 : nand02 port map ( Y=>nx14093, A0=>nx35783, A1=>nx25832);
   ix13834 : mux21_ni port map ( Y=>nx13833, A0=>num_in_2, A1=>num_out_2, S0
      =>nx35795);
   ix497 : ao22 port map ( Y=>nx496, A0=>mdr_data_out(2), A1=>nx12893, B0=>
      nx35625, B1=>nx35713);
   ix35624 : inv01 port map ( Y=>nx35625, A=>nx25821);
   ix13664 : mux21 port map ( Y=>nx13663, A0=>nx35153, A1=>nx35799, S0=>
      nx35097);
   ix13714 : mux21_ni port map ( Y=>nx13713, A0=>num_in_0, A1=>num_out_0, S0
      =>nx35795);
   ix377 : ao22 port map ( Y=>nx376, A0=>mdr_data_out(0), A1=>nx12893, B0=>
      nx35627, B1=>nx35713);
   ix35626 : inv01 port map ( Y=>nx35627, A=>nx25864);
   ix805 : and03 port map ( Y=>nx12879, A0=>nx25857, A1=>nx35783, A2=>
      state(1));
   ix173 : and03 port map ( Y=>nx172, A0=>state(0), A1=>nx35783, A2=>nx35779
   );
   ix25860 : nor03_2x port map ( Y=>nx4, A0=>nx25857, A1=>state(2), A2=>
      nx35779);
   ix811 : ao21 port map ( Y=>nx12877, A0=>nx25857, A1=>nx35779, B0=>nx35783
   );
   ix25865 : xor2 port map ( Y=>nx25864, A0=>alu_inp1_0, A1=>nx25935);
   ix391 : mux21_ni port map ( Y=>nx390, A0=>address_out_0, A1=>num_out_0, 
      S0=>nx35713);
   ix25875 : nor02ii port map ( Y=>nx25874, A0=>sub_state(1), A1=>nx12893);
   ix27 : nor02ii port map ( Y=>nx26, A0=>nx25879, A1=>nx12887);
   ix21 : ao32 port map ( Y=>nx20, A0=>nx12887, A1=>nx35791, A2=>nx35629, B0
      =>nx25944, B1=>nx35713);
   ix35628 : inv01 port map ( Y=>nx35629, A=>nx34401);
   ix175 : and02 port map ( Y=>nx174, A0=>nx35785, A1=>nx35779);
   ix25890 : nand02 port map ( Y=>nx12882, A0=>nx35915, A1=>nx35589);
   ix25894 : nor02ii port map ( Y=>nx25893, A0=>nx174, A1=>nx35153);
   ix335 : ao32 port map ( Y=>nx334, A0=>nx35631, A1=>nx35791, A2=>nx320, B0
      =>nx35101, B1=>nx25907);
   ix25906 : nand02 port map ( Y=>nx35631, A0=>nx186, A1=>nx172);
   ix25908 : nor02ii port map ( Y=>nx25907, A0=>nx35157, A1=>nx35791);
   ix225 : and03 port map ( Y=>nx12893, A0=>nx25857, A1=>nx35785, A2=>
      nx35781);
   ix243 : mux21 port map ( Y=>nx242, A0=>nx35793, A1=>nx35153, S0=>nx35101
   );
   ix13774 : mux21_ni port map ( Y=>nx13773, A0=>num_in_1, A1=>num_out_1, S0
      =>nx35795);
   ix413 : mux21_ni port map ( Y=>nx412, A0=>alu_inp1_0, A1=>nx34499, S0=>
      nx25935);
   ix25963 : xor2 port map ( Y=>nx25962, A0=>alu_inp1_1, A1=>nx35799);
   ix449 : mux21_ni port map ( Y=>nx448, A0=>address_out_1, A1=>num_out_1, 
      S0=>nx35713);
   ix13884 : mux21_ni port map ( Y=>nx13883, A0=>num_in_3, A1=>num_out_3, S0
      =>nx35795);
   ix25987 : xnor2 port map ( Y=>nx25986, A0=>nx25998, A1=>nx35799);
   ix481 : mux21_ni port map ( Y=>nx480, A0=>address_out_2, A1=>num_out_2, 
      S0=>nx35715);
   ix26002 : xor2 port map ( Y=>nx26001, A0=>alu_inp1_3, A1=>nx35801);
   ix541 : mux21_ni port map ( Y=>nx540, A0=>address_out_3, A1=>num_out_3, 
      S0=>nx35715);
   ix13934 : mux21_ni port map ( Y=>nx13933, A0=>num_in_4, A1=>num_out_4, S0
      =>nx35795);
   ix607 : ao22 port map ( Y=>nx606, A0=>mdr_data_out(4), A1=>nx12893, B0=>
      nx35633, B1=>nx35715);
   ix35632 : inv01 port map ( Y=>nx35633, A=>nx26022);
   ix26028 : xnor2 port map ( Y=>nx26027, A0=>nx26039, A1=>nx35801);
   ix591 : mux21_ni port map ( Y=>nx590, A0=>address_out_4, A1=>num_out_4, 
      S0=>nx35715);
   ix26045 : or04 port map ( Y=>nx26044, A0=>num_out_5, A1=>num_out_6, A2=>
      num_out_7, A3=>nx35917);
   ix13984 : mux21 port map ( Y=>nx13983, A0=>nx26069, A1=>nx26046, S0=>
      nx35795);
   ix26057 : xor2 port map ( Y=>nx26056, A0=>alu_inp1_5, A1=>nx35801);
   ix649 : mux21_ni port map ( Y=>nx648, A0=>address_out_5, A1=>num_out_5, 
      S0=>nx35715);
   ix14034 : mux21_ni port map ( Y=>nx14033, A0=>num_in_6, A1=>num_out_6, S0
      =>nx35797);
   ix715 : ao22 port map ( Y=>nx714, A0=>mdr_data_out(6), A1=>nx12893, B0=>
      nx35635, B1=>nx35715);
   ix35634 : inv01 port map ( Y=>nx35635, A=>nx26078);
   ix26084 : xnor2 port map ( Y=>nx26083, A0=>nx26095, A1=>nx35801);
   ix699 : mux21_ni port map ( Y=>nx698, A0=>address_out_6, A1=>num_out_6, 
      S0=>nx35715);
   ix14084 : mux21 port map ( Y=>nx14083, A0=>nx26122, A1=>nx26099, S0=>
      nx35797);
   ix26110 : xor2 port map ( Y=>nx26109, A0=>alu_inp1_7, A1=>nx35801);
   ix755 : mux21_ni port map ( Y=>nx754, A0=>address_out_7, A1=>num_out_7, 
      S0=>nx35717);
   ix843 : and03 port map ( Y=>nx12909, A0=>nx25857, A1=>state(2), A2=>
      nx35781);
   ix26140 : oai21 port map ( Y=>nx35621, A0=>nx35793, A1=>nx35101, B0=>
      nx35637);
   ix819 : or04 port map ( Y=>nx35637, A0=>nx12891, A1=>nx25900, A2=>nx35155, 
      A3=>nx35157);
   ix65 : and04 port map ( Y=>nx64, A0=>nx35785, A1=>state(1), A2=>nx35639, 
      A3=>nx25942);
   ix35638 : inv01 port map ( Y=>nx35639, A=>nx56);
   ix26183 : or02 port map ( Y=>nx26182, A0=>nx26176, A1=>max_calc_start);
   ix26192 : and02 port map ( Y=>nx26191, A0=>nx26176, A1=>nx26180);
   ix26195 : xnor2 port map ( Y=>nx26194, A0=>nx26188, A1=>nx35977);
   ix17554 : ao32 port map ( Y=>nx17553, A0=>nx35641, A1=>nx26203, A2=>
      max_calc_start, B0=>nx36331, B1=>nx26191);
   ix35640 : inv01 port map ( Y=>nx35641, A=>nx26194);
   ix17564 : ao22 port map ( Y=>nx17563, A0=>max_calc_start, A1=>nx35843, B0
      =>max_calc_state_3, B1=>nx26191);
   ix6277 : nor03_2x port map ( Y=>nx34735, A0=>nx26188, A1=>nx35977, A2=>
      nx35643);
   ix35642 : inv01 port map ( Y=>nx35643, A=>nx26201);
   ix26202 : and02 port map ( Y=>nx26201, A0=>nx36299, A1=>nx26203);
   ix25564 : mux21_ni port map ( Y=>nx25563, A0=>answer_0_EXMPLR, A1=>
      nx13121, S0=>nx35741);
   ix19151 : mux21_ni port map ( Y=>nx13121, A0=>
      max_calc_comparator_first_inp2_0, A1=>max_calc_comparator_first_inp1_0, 
      S0=>nx35905);
   ix19634 : mux21_ni port map ( Y=>nx19633, A0=>
      max_calc_comparator_first_inp1_0, A1=>nx9512, S0=>nx36281);
   ix9513 : mux21_ni port map ( Y=>nx9512, A0=>nx9508, A1=>nx6388, S0=>
      nx35959);
   ix6389 : mux21_ni port map ( Y=>nx6388, A0=>max_calc_ans1_0, A1=>
      label_1_output(0), S0=>nx35977);
   ix17224 : mux21_ni port map ( Y=>nx17223, A0=>label_1_output(0), A1=>
      label_1_input_0, S0=>nx36241);
   ix17214 : mux21_ni port map ( Y=>nx17213, A0=>
      label_1_input_state_machine_0, A1=>mdr_data_out(0), S0=>nx36201);
   ix17204 : mux21_ni port map ( Y=>nx17203, A0=>nx35731, A1=>nx5736, S0=>
      nx35199);
   ix5737 : mux21_ni port map ( Y=>nx5736, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_0_1, S0=>nx36011);
   ix17194 : mux21_ni port map ( Y=>nx17193, A0=>
      booth_booth_integration_output_0_1, A1=>nx5724, S0=>nx35199);
   ix5725 : mux21_ni port map ( Y=>nx5724, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_0_2, S0=>nx36011);
   ix17184 : mux21_ni port map ( Y=>nx17183, A0=>
      booth_booth_integration_output_0_2, A1=>nx5712, S0=>nx35199);
   ix5713 : mux21_ni port map ( Y=>nx5712, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_0_3, S0=>nx36011);
   ix17174 : mux21_ni port map ( Y=>nx17173, A0=>
      booth_booth_integration_output_0_3, A1=>nx5700, S0=>nx35199);
   ix5701 : mux21_ni port map ( Y=>nx5700, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_0_4, S0=>nx36011);
   ix17164 : mux21_ni port map ( Y=>nx17163, A0=>
      booth_booth_integration_output_0_4, A1=>nx5688, S0=>nx35199);
   ix5689 : mux21_ni port map ( Y=>nx5688, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_0_5, S0=>nx36011);
   ix17154 : mux21_ni port map ( Y=>nx17153, A0=>
      booth_booth_integration_output_0_5, A1=>nx5676, S0=>nx35199);
   ix5677 : mux21_ni port map ( Y=>nx5676, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_0_6, S0=>nx36013);
   ix17144 : mux21_ni port map ( Y=>nx17143, A0=>
      booth_booth_integration_output_0_6, A1=>nx5664, S0=>nx35199);
   ix5665 : mux21_ni port map ( Y=>nx5664, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_0_7, S0=>nx36013);
   ix17134 : mux21_ni port map ( Y=>nx17133, A0=>
      booth_booth_integration_output_0_7, A1=>nx5652, S0=>nx36003);
   ix5653 : mux21_ni port map ( Y=>nx5652, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_0_8, S0=>nx36013);
   ix17124 : mux21_ni port map ( Y=>nx17123, A0=>
      booth_booth_integration_output_0_8, A1=>nx5640, S0=>nx36003);
   ix5641 : mux21_ni port map ( Y=>nx5640, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_0_9, S0=>nx36013);
   ix17114 : mux21_ni port map ( Y=>nx17113, A0=>
      booth_booth_integration_output_0_9, A1=>nx5628, S0=>nx36003);
   ix5629 : mux21_ni port map ( Y=>nx5628, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_0_10, S0=>nx36013);
   ix17104 : mux21_ni port map ( Y=>nx17103, A0=>
      booth_booth_integration_output_0_10, A1=>nx5616, S0=>nx36005);
   ix5617 : mux21_ni port map ( Y=>nx5616, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_0_11, S0=>nx36013);
   ix17094 : mux21_ni port map ( Y=>nx17093, A0=>
      booth_booth_integration_output_0_11, A1=>nx5604, S0=>nx36005);
   ix5605 : mux21_ni port map ( Y=>nx5604, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_0_12, S0=>nx36013);
   ix17084 : mux21_ni port map ( Y=>nx17083, A0=>
      booth_booth_integration_output_0_12, A1=>nx5592, S0=>nx36005);
   ix5593 : mux21_ni port map ( Y=>nx5592, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_0_13, S0=>nx36015);
   ix17074 : mux21_ni port map ( Y=>nx17073, A0=>
      booth_booth_integration_output_0_13, A1=>nx5580, S0=>nx36005);
   ix5581 : mux21_ni port map ( Y=>nx5580, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_0_14, S0=>nx36015);
   ix17064 : mux21_ni port map ( Y=>nx17063, A0=>
      booth_booth_integration_output_0_14, A1=>nx5568, S0=>nx36005);
   ix5569 : mux21_ni port map ( Y=>nx5568, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_0_15, S0=>nx36015);
   ix17054 : mux21 port map ( Y=>nx17053, A0=>nx26634, A1=>nx26276, S0=>
      nx36005);
   ix16704 : mux21_ni port map ( Y=>nx16703, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_0, A1=>nx34667, S0=>nx35803
   );
   ix16690 : and02 port map ( Y=>nx16689, A0=>nx36327, A1=>
      booth_booth_integrtaion_0_shift_Reg_count_0);
   ix16884 : mux21_ni port map ( Y=>nx16883, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_9, A1=>nx34653, S0=>nx35803
   );
   ix16874 : mux21_ni port map ( Y=>nx16873, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_8, S0=>nx36005);
   ix16864 : mux21_ni port map ( Y=>nx16863, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_8, S0=>nx35803);
   ix16854 : mux21_ni port map ( Y=>nx16853, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_7, S0=>nx36007);
   ix16844 : mux21_ni port map ( Y=>nx16843, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_7, S0=>nx35803);
   ix16834 : mux21_ni port map ( Y=>nx16833, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_6, S0=>nx36007);
   ix16824 : mux21_ni port map ( Y=>nx16823, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_6, S0=>nx35803);
   ix16814 : mux21_ni port map ( Y=>nx16813, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_5, S0=>nx36007);
   ix16804 : mux21_ni port map ( Y=>nx16803, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_5, S0=>nx35803);
   ix16794 : mux21_ni port map ( Y=>nx16793, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_4, S0=>nx36007);
   ix16784 : mux21_ni port map ( Y=>nx16783, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_4, S0=>nx35805);
   ix16774 : mux21_ni port map ( Y=>nx16773, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_3, S0=>nx36007);
   ix16764 : mux21_ni port map ( Y=>nx16763, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_3, S0=>nx35805);
   ix16754 : mux21_ni port map ( Y=>nx16753, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_2, S0=>nx36007);
   ix16744 : mux21_ni port map ( Y=>nx16743, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_2, S0=>nx35805);
   ix16734 : mux21_ni port map ( Y=>nx16733, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_1, S0=>nx36007);
   ix16724 : mux21_ni port map ( Y=>nx16723, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_0_shift_Reg_output_1, S0=>nx35805);
   ix16714 : mux21_ni port map ( Y=>nx16713, A0=>
      booth_booth_integrtaion_0_shift_Reg_count_1, A1=>nx34667, S0=>nx36009
   );
   ix5009 : and02 port map ( Y=>nx5008, A0=>nx26349, A1=>nx35731);
   ix26352 : or03 port map ( Y=>nx26351, A0=>nx26353, A1=>
      booth_booth_integrtaion_0_shift_reg_output_0, A2=>nx36327);
   ix17044 : mux21_ni port map ( Y=>nx17043, A0=>
      booth_booth_integrtaion_0_booth_output_16, A1=>nx5538, S0=>nx36009);
   ix5539 : nor02ii port map ( Y=>nx5538, A0=>nx26360, A1=>nx36015);
   ix5015 : nor02ii port map ( Y=>nx5014, A0=>nx26344, A1=>
      booth_booth_integrtaion_0_booth_output_16);
   ix5533 : xor2 port map ( Y=>nx13067, A0=>nx26366, A1=>nx26630);
   ix5521 : xor2 port map ( Y=>nx13069, A0=>nx26391, A1=>nx35205);
   ix17024 : mux21_ni port map ( Y=>nx17023, A0=>
      booth_booth_integrtaion_0_booth_output_18, A1=>nx5514, S0=>nx36009);
   ix5515 : nor02ii port map ( Y=>nx5514, A0=>nx26381, A1=>nx36015);
   ix5509 : xor2 port map ( Y=>nx13071, A0=>nx26396, A1=>nx26627);
   ix26413 : or02 port map ( Y=>nx26412, A0=>nx26349, A1=>nx35733);
   ix5497 : xor2 port map ( Y=>nx13073, A0=>nx26430, A1=>nx35207);
   ix17004 : mux21_ni port map ( Y=>nx17003, A0=>
      booth_booth_integrtaion_0_booth_output_20, A1=>nx5490, S0=>nx36009);
   ix5491 : nor02ii port map ( Y=>nx5490, A0=>nx26418, A1=>nx36015);
   ix5485 : xor2 port map ( Y=>nx13074, A0=>nx26435, A1=>nx26624);
   ix5473 : xor2 port map ( Y=>nx13075, A0=>nx26465, A1=>nx35209);
   ix16984 : mux21_ni port map ( Y=>nx16983, A0=>
      booth_booth_integrtaion_0_booth_output_22, A1=>nx5466, S0=>nx36009);
   ix5467 : nor02ii port map ( Y=>nx5466, A0=>nx26453, A1=>nx36015);
   ix5461 : xor2 port map ( Y=>nx13077, A0=>nx26470, A1=>nx26621);
   ix5449 : xor2 port map ( Y=>nx13079, A0=>nx26500, A1=>nx35211);
   ix16964 : mux21_ni port map ( Y=>nx16963, A0=>
      booth_booth_integrtaion_0_booth_output_24, A1=>nx5442, S0=>nx36009);
   ix5443 : nor02ii port map ( Y=>nx5442, A0=>nx26488, A1=>nx36017);
   ix5437 : xor2 port map ( Y=>nx13081, A0=>nx26505, A1=>nx26618);
   ix5425 : xor2 port map ( Y=>nx13083, A0=>nx26535, A1=>nx35213);
   ix16944 : mux21_ni port map ( Y=>nx16943, A0=>
      booth_booth_integrtaion_0_booth_output_26, A1=>nx5418, S0=>nx36009);
   ix5419 : nor02ii port map ( Y=>nx5418, A0=>nx26523, A1=>nx36017);
   ix5413 : xor2 port map ( Y=>nx13085, A0=>nx26540, A1=>nx26615);
   ix5401 : xor2 port map ( Y=>nx13087, A0=>nx26570, A1=>nx35215);
   ix16924 : mux21_ni port map ( Y=>nx16923, A0=>
      booth_booth_integrtaion_0_booth_output_28, A1=>nx5394, S0=>nx35197);
   ix5395 : nor02ii port map ( Y=>nx5394, A0=>nx26558, A1=>nx36017);
   ix5389 : xor2 port map ( Y=>nx13089, A0=>nx26575, A1=>nx26612);
   ix5377 : xor2 port map ( Y=>nx13090, A0=>nx26605, A1=>nx35217);
   ix16904 : mux21_ni port map ( Y=>nx16903, A0=>
      booth_booth_integrtaion_0_booth_output_31, A1=>nx5370, S0=>nx35197);
   ix5371 : nor02ii port map ( Y=>nx5370, A0=>nx26593, A1=>nx36017);
   ix5365 : xor2 port map ( Y=>nx5364, A0=>nx26605, A1=>nx26608);
   ix5551 : nor02ii port map ( Y=>nx5550, A0=>nx5014, A1=>nx36017);
   ix26658 : oai21 port map ( Y=>nx846, A0=>nx35781, A1=>nx25857, B0=>
      nx35785);
   ix26667 : and02 port map ( Y=>nx26666, A0=>nx35791, A1=>sub_state(1));
   ix26670 : nor02ii port map ( Y=>nx26669, A0=>sel_dst_0, A1=>nx35919);
   ix17584 : mux21_ni port map ( Y=>nx17583, A0=>nx13121, A1=>
      max_calc_ans1_0, S0=>nx35851);
   ix6379 : nand03 port map ( Y=>nx34821, A0=>nx35959, A1=>nx26203, A2=>
      nx36291);
   ix9509 : mux21_ni port map ( Y=>nx9508, A0=>max_calc_ans5_0, A1=>
      max_calc_ans6_0, S0=>nx35977);
   ix17594 : mux21_ni port map ( Y=>nx17593, A0=>max_calc_ans6_0, A1=>
      nx13121, S0=>nx36021);
   ix26683 : nor02ii port map ( Y=>nx35289, A0=>nx36381, A1=>nx26194);
   ix19624 : mux21_ni port map ( Y=>nx19623, A0=>max_calc_ans5_0, A1=>nx9498, 
      S0=>nx36291);
   ix9499 : mux21 port map ( Y=>nx9498, A0=>nx27133, A1=>nx26693, S0=>
      nx35861);
   ix18144 : mux21_ni port map ( Y=>nx18143, A0=>label_9_output(0), A1=>
      label_9_input_0, S0=>nx36241);
   ix18134 : mux21_ni port map ( Y=>nx18133, A0=>
      label_9_input_state_machine_0, A1=>mdr_data_out(128), S0=>nx36201);
   ix18124 : mux21_ni port map ( Y=>nx18123, A0=>nx35755, A1=>nx7236, S0=>
      nx35307);
   ix7237 : mux21_ni port map ( Y=>nx7236, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_8_1, S0=>nx36039);
   ix18114 : mux21_ni port map ( Y=>nx18113, A0=>
      booth_booth_integration_output_8_1, A1=>nx7224, S0=>nx35307);
   ix7225 : mux21_ni port map ( Y=>nx7224, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_8_2, S0=>nx36039);
   ix18104 : mux21_ni port map ( Y=>nx18103, A0=>
      booth_booth_integration_output_8_2, A1=>nx7212, S0=>nx35307);
   ix7213 : mux21_ni port map ( Y=>nx7212, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_8_3, S0=>nx36039);
   ix18094 : mux21_ni port map ( Y=>nx18093, A0=>
      booth_booth_integration_output_8_3, A1=>nx7200, S0=>nx35307);
   ix7201 : mux21_ni port map ( Y=>nx7200, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_8_4, S0=>nx36039);
   ix18084 : mux21_ni port map ( Y=>nx18083, A0=>
      booth_booth_integration_output_8_4, A1=>nx7188, S0=>nx35307);
   ix7189 : mux21_ni port map ( Y=>nx7188, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_8_5, S0=>nx36039);
   ix18074 : mux21_ni port map ( Y=>nx18073, A0=>
      booth_booth_integration_output_8_5, A1=>nx7176, S0=>nx35307);
   ix7177 : mux21_ni port map ( Y=>nx7176, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_8_6, S0=>nx36041);
   ix18064 : mux21_ni port map ( Y=>nx18063, A0=>
      booth_booth_integration_output_8_6, A1=>nx7164, S0=>nx35307);
   ix7165 : mux21_ni port map ( Y=>nx7164, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_8_7, S0=>nx36041);
   ix18054 : mux21_ni port map ( Y=>nx18053, A0=>
      booth_booth_integration_output_8_7, A1=>nx7152, S0=>nx36031);
   ix7153 : mux21_ni port map ( Y=>nx7152, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_8_8, S0=>nx36041);
   ix18044 : mux21_ni port map ( Y=>nx18043, A0=>
      booth_booth_integration_output_8_8, A1=>nx7140, S0=>nx36031);
   ix7141 : mux21_ni port map ( Y=>nx7140, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_8_9, S0=>nx36041);
   ix18034 : mux21_ni port map ( Y=>nx18033, A0=>
      booth_booth_integration_output_8_9, A1=>nx7128, S0=>nx36031);
   ix7129 : mux21_ni port map ( Y=>nx7128, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_8_10, S0=>nx36041);
   ix18024 : mux21_ni port map ( Y=>nx18023, A0=>
      booth_booth_integration_output_8_10, A1=>nx7116, S0=>nx36033);
   ix7117 : mux21_ni port map ( Y=>nx7116, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_8_11, S0=>nx36041);
   ix18014 : mux21_ni port map ( Y=>nx18013, A0=>
      booth_booth_integration_output_8_11, A1=>nx7104, S0=>nx36033);
   ix7105 : mux21_ni port map ( Y=>nx7104, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_8_12, S0=>nx36041);
   ix18004 : mux21_ni port map ( Y=>nx18003, A0=>
      booth_booth_integration_output_8_12, A1=>nx7092, S0=>nx36033);
   ix7093 : mux21_ni port map ( Y=>nx7092, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_8_13, S0=>nx36043);
   ix17994 : mux21_ni port map ( Y=>nx17993, A0=>
      booth_booth_integration_output_8_13, A1=>nx7080, S0=>nx36033);
   ix7081 : mux21_ni port map ( Y=>nx7080, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_8_14, S0=>nx36043);
   ix17984 : mux21_ni port map ( Y=>nx17983, A0=>
      booth_booth_integration_output_8_14, A1=>nx7068, S0=>nx36033);
   ix7069 : mux21_ni port map ( Y=>nx7068, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_8_15, S0=>nx36043);
   ix17974 : mux21 port map ( Y=>nx17973, A0=>nx27113, A1=>nx26755, S0=>
      nx36033);
   ix17624 : mux21_ni port map ( Y=>nx17623, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_0, A1=>nx34847, S0=>nx35807
   );
   ix17610 : and02 port map ( Y=>nx17609, A0=>nx36341, A1=>
      booth_booth_integrtaion_8_shift_Reg_count_0);
   ix17804 : mux21_ni port map ( Y=>nx17803, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_9, A1=>nx34833, S0=>nx35807
   );
   ix17794 : mux21_ni port map ( Y=>nx17793, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_8, S0=>nx36033);
   ix17784 : mux21_ni port map ( Y=>nx17783, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_8, S0=>nx35807);
   ix17774 : mux21_ni port map ( Y=>nx17773, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_7, S0=>nx36035);
   ix17764 : mux21_ni port map ( Y=>nx17763, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_7, S0=>nx35807);
   ix17754 : mux21_ni port map ( Y=>nx17753, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_6, S0=>nx36035);
   ix17744 : mux21_ni port map ( Y=>nx17743, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_6, S0=>nx35807);
   ix17734 : mux21_ni port map ( Y=>nx17733, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_5, S0=>nx36035);
   ix17724 : mux21_ni port map ( Y=>nx17723, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_5, S0=>nx35807);
   ix17714 : mux21_ni port map ( Y=>nx17713, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_4, S0=>nx36035);
   ix17704 : mux21_ni port map ( Y=>nx17703, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_4, S0=>nx35809);
   ix17694 : mux21_ni port map ( Y=>nx17693, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_3, S0=>nx36035);
   ix17684 : mux21_ni port map ( Y=>nx17683, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_3, S0=>nx35809);
   ix17674 : mux21_ni port map ( Y=>nx17673, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_2, S0=>nx36035);
   ix17664 : mux21_ni port map ( Y=>nx17663, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_2, S0=>nx35809);
   ix17654 : mux21_ni port map ( Y=>nx17653, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_1, S0=>nx36035);
   ix17644 : mux21_ni port map ( Y=>nx17643, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_8_shift_Reg_output_1, S0=>nx35809);
   ix17634 : mux21_ni port map ( Y=>nx17633, A0=>
      booth_booth_integrtaion_8_shift_Reg_count_1, A1=>nx34847, S0=>nx36037
   );
   ix6509 : and02 port map ( Y=>nx6508, A0=>nx26828, A1=>nx35755);
   ix26831 : or03 port map ( Y=>nx26830, A0=>nx26832, A1=>
      booth_booth_integrtaion_8_shift_reg_output_0, A2=>nx36341);
   ix17964 : mux21_ni port map ( Y=>nx17963, A0=>
      booth_booth_integrtaion_8_booth_output_16, A1=>nx7038, S0=>nx36037);
   ix7039 : nor02ii port map ( Y=>nx7038, A0=>nx26839, A1=>nx36043);
   ix6515 : nor02ii port map ( Y=>nx6514, A0=>nx26823, A1=>
      booth_booth_integrtaion_8_booth_output_16);
   ix7033 : xor2 port map ( Y=>nx13123, A0=>nx26845, A1=>nx27109);
   ix7021 : xor2 port map ( Y=>nx13125, A0=>nx26870, A1=>nx35313);
   ix17944 : mux21_ni port map ( Y=>nx17943, A0=>
      booth_booth_integrtaion_8_booth_output_18, A1=>nx7014, S0=>nx36037);
   ix7015 : nor02ii port map ( Y=>nx7014, A0=>nx26860, A1=>nx36043);
   ix7009 : xor2 port map ( Y=>nx13127, A0=>nx26875, A1=>nx27106);
   ix26892 : or02 port map ( Y=>nx26891, A0=>nx26828, A1=>nx35757);
   ix6997 : xor2 port map ( Y=>nx13129, A0=>nx26909, A1=>nx35315);
   ix17924 : mux21_ni port map ( Y=>nx17923, A0=>
      booth_booth_integrtaion_8_booth_output_20, A1=>nx6990, S0=>nx36037);
   ix6991 : nor02ii port map ( Y=>nx6990, A0=>nx26897, A1=>nx36043);
   ix6985 : xor2 port map ( Y=>nx13131, A0=>nx26914, A1=>nx27103);
   ix6973 : xor2 port map ( Y=>nx13133, A0=>nx26944, A1=>nx35317);
   ix17904 : mux21_ni port map ( Y=>nx17903, A0=>
      booth_booth_integrtaion_8_booth_output_22, A1=>nx6966, S0=>nx36037);
   ix6967 : nor02ii port map ( Y=>nx6966, A0=>nx26932, A1=>nx36043);
   ix6961 : xor2 port map ( Y=>nx13135, A0=>nx26949, A1=>nx27100);
   ix6949 : xor2 port map ( Y=>nx13137, A0=>nx26979, A1=>nx35319);
   ix17884 : mux21_ni port map ( Y=>nx17883, A0=>
      booth_booth_integrtaion_8_booth_output_24, A1=>nx6942, S0=>nx36037);
   ix6943 : nor02ii port map ( Y=>nx6942, A0=>nx26967, A1=>nx36045);
   ix6937 : xor2 port map ( Y=>nx13138, A0=>nx26984, A1=>nx27097);
   ix6925 : xor2 port map ( Y=>nx13139, A0=>nx27014, A1=>nx35321);
   ix17864 : mux21_ni port map ( Y=>nx17863, A0=>
      booth_booth_integrtaion_8_booth_output_26, A1=>nx6918, S0=>nx36037);
   ix6919 : nor02ii port map ( Y=>nx6918, A0=>nx27002, A1=>nx36045);
   ix6913 : xor2 port map ( Y=>nx13141, A0=>nx27019, A1=>nx27094);
   ix6901 : xor2 port map ( Y=>nx13143, A0=>nx27049, A1=>nx35323);
   ix17844 : mux21_ni port map ( Y=>nx17843, A0=>
      booth_booth_integrtaion_8_booth_output_28, A1=>nx6894, S0=>nx35305);
   ix6895 : nor02ii port map ( Y=>nx6894, A0=>nx27037, A1=>nx36045);
   ix6889 : xor2 port map ( Y=>nx13145, A0=>nx27054, A1=>nx27091);
   ix6877 : xor2 port map ( Y=>nx13146, A0=>nx27084, A1=>nx35325);
   ix17824 : mux21_ni port map ( Y=>nx17823, A0=>
      booth_booth_integrtaion_8_booth_output_31, A1=>nx6870, S0=>nx35305);
   ix6871 : nor02ii port map ( Y=>nx6870, A0=>nx27072, A1=>nx36045);
   ix6865 : xor2 port map ( Y=>nx6864, A0=>nx27084, A1=>nx27087);
   ix7051 : nor02ii port map ( Y=>nx7050, A0=>nx6514, A1=>nx36045);
   ix18714 : mux21_ni port map ( Y=>nx18713, A0=>label_10_output(0), A1=>
      label_10_input_0, S0=>nx36241);
   ix18704 : mux21_ni port map ( Y=>nx18703, A0=>
      label_10_input_state_machine_0, A1=>mdr_data_out(144), S0=>nx36201);
   ix18694 : mux21_ni port map ( Y=>nx18693, A0=>nx35759, A1=>nx8116, S0=>
      nx35333);
   ix8117 : mux21_ni port map ( Y=>nx8116, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_9_1, S0=>nx36055);
   ix18684 : mux21_ni port map ( Y=>nx18683, A0=>
      booth_booth_integration_output_9_1, A1=>nx8104, S0=>nx35333);
   ix8105 : mux21_ni port map ( Y=>nx8104, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_9_2, S0=>nx36055);
   ix18674 : mux21_ni port map ( Y=>nx18673, A0=>
      booth_booth_integration_output_9_2, A1=>nx8092, S0=>nx35333);
   ix8093 : mux21_ni port map ( Y=>nx8092, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_9_3, S0=>nx36055);
   ix18664 : mux21_ni port map ( Y=>nx18663, A0=>
      booth_booth_integration_output_9_3, A1=>nx8080, S0=>nx35333);
   ix8081 : mux21_ni port map ( Y=>nx8080, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_9_4, S0=>nx36055);
   ix18654 : mux21_ni port map ( Y=>nx18653, A0=>
      booth_booth_integration_output_9_4, A1=>nx8068, S0=>nx35333);
   ix8069 : mux21_ni port map ( Y=>nx8068, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_9_5, S0=>nx36055);
   ix18644 : mux21_ni port map ( Y=>nx18643, A0=>
      booth_booth_integration_output_9_5, A1=>nx8056, S0=>nx35333);
   ix8057 : mux21_ni port map ( Y=>nx8056, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_9_6, S0=>nx36057);
   ix18634 : mux21_ni port map ( Y=>nx18633, A0=>
      booth_booth_integration_output_9_6, A1=>nx8044, S0=>nx35333);
   ix8045 : mux21_ni port map ( Y=>nx8044, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_9_7, S0=>nx36057);
   ix18624 : mux21_ni port map ( Y=>nx18623, A0=>
      booth_booth_integration_output_9_7, A1=>nx8032, S0=>nx36047);
   ix8033 : mux21_ni port map ( Y=>nx8032, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_9_8, S0=>nx36057);
   ix18614 : mux21_ni port map ( Y=>nx18613, A0=>
      booth_booth_integration_output_9_8, A1=>nx8020, S0=>nx36047);
   ix8021 : mux21_ni port map ( Y=>nx8020, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_9_9, S0=>nx36057);
   ix18604 : mux21_ni port map ( Y=>nx18603, A0=>
      booth_booth_integration_output_9_9, A1=>nx8008, S0=>nx36047);
   ix8009 : mux21_ni port map ( Y=>nx8008, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_9_10, S0=>nx36057);
   ix18594 : mux21_ni port map ( Y=>nx18593, A0=>
      booth_booth_integration_output_9_10, A1=>nx7996, S0=>nx36049);
   ix7997 : mux21_ni port map ( Y=>nx7996, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_9_11, S0=>nx36057);
   ix18584 : mux21_ni port map ( Y=>nx18583, A0=>
      booth_booth_integration_output_9_11, A1=>nx7984, S0=>nx36049);
   ix7985 : mux21_ni port map ( Y=>nx7984, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_9_12, S0=>nx36057);
   ix18574 : mux21_ni port map ( Y=>nx18573, A0=>
      booth_booth_integration_output_9_12, A1=>nx7972, S0=>nx36049);
   ix7973 : mux21_ni port map ( Y=>nx7972, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_9_13, S0=>nx36059);
   ix18564 : mux21_ni port map ( Y=>nx18563, A0=>
      booth_booth_integration_output_9_13, A1=>nx7960, S0=>nx36049);
   ix7961 : mux21_ni port map ( Y=>nx7960, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_9_14, S0=>nx36059);
   ix18554 : mux21_ni port map ( Y=>nx18553, A0=>
      booth_booth_integration_output_9_14, A1=>nx7948, S0=>nx36049);
   ix7949 : mux21_ni port map ( Y=>nx7948, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_9_15, S0=>nx36059);
   ix18544 : mux21 port map ( Y=>nx18543, A0=>nx27552, A1=>nx27194, S0=>
      nx36049);
   ix18194 : mux21_ni port map ( Y=>nx18193, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_0, A1=>nx34879, S0=>nx35811
   );
   ix18180 : and02 port map ( Y=>nx18179, A0=>nx36345, A1=>
      booth_booth_integrtaion_9_shift_Reg_count_0);
   ix18374 : mux21_ni port map ( Y=>nx18373, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_9, A1=>nx34865, S0=>nx35811
   );
   ix18364 : mux21_ni port map ( Y=>nx18363, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_8, S0=>nx36049);
   ix18354 : mux21_ni port map ( Y=>nx18353, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_8, S0=>nx35811);
   ix18344 : mux21_ni port map ( Y=>nx18343, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_7, S0=>nx36051);
   ix18334 : mux21_ni port map ( Y=>nx18333, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_7, S0=>nx35811);
   ix18324 : mux21_ni port map ( Y=>nx18323, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_6, S0=>nx36051);
   ix18314 : mux21_ni port map ( Y=>nx18313, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_6, S0=>nx35811);
   ix18304 : mux21_ni port map ( Y=>nx18303, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_5, S0=>nx36051);
   ix18294 : mux21_ni port map ( Y=>nx18293, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_5, S0=>nx35811);
   ix18284 : mux21_ni port map ( Y=>nx18283, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_4, S0=>nx36051);
   ix18274 : mux21_ni port map ( Y=>nx18273, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_4, S0=>nx35813);
   ix18264 : mux21_ni port map ( Y=>nx18263, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_3, S0=>nx36051);
   ix18254 : mux21_ni port map ( Y=>nx18253, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_3, S0=>nx35813);
   ix18244 : mux21_ni port map ( Y=>nx18243, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_2, S0=>nx36051);
   ix18234 : mux21_ni port map ( Y=>nx18233, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_2, S0=>nx35813);
   ix18224 : mux21_ni port map ( Y=>nx18223, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_1, S0=>nx36051);
   ix18214 : mux21_ni port map ( Y=>nx18213, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_9_shift_Reg_output_1, S0=>nx35813);
   ix18204 : mux21_ni port map ( Y=>nx18203, A0=>
      booth_booth_integrtaion_9_shift_Reg_count_1, A1=>nx34879, S0=>nx36053
   );
   ix7389 : and02 port map ( Y=>nx7388, A0=>nx27267, A1=>nx35759);
   ix27270 : or03 port map ( Y=>nx27269, A0=>nx27271, A1=>
      booth_booth_integrtaion_9_shift_reg_output_0, A2=>nx36345);
   ix18534 : mux21_ni port map ( Y=>nx18533, A0=>
      booth_booth_integrtaion_9_booth_output_16, A1=>nx7918, S0=>nx36053);
   ix7919 : nor02ii port map ( Y=>nx7918, A0=>nx27278, A1=>nx36059);
   ix7395 : nor02ii port map ( Y=>nx7394, A0=>nx27262, A1=>
      booth_booth_integrtaion_9_booth_output_16);
   ix7913 : xor2 port map ( Y=>nx13149, A0=>nx27284, A1=>nx27548);
   ix7901 : xor2 port map ( Y=>nx13151, A0=>nx27309, A1=>nx35339);
   ix18514 : mux21_ni port map ( Y=>nx18513, A0=>
      booth_booth_integrtaion_9_booth_output_18, A1=>nx7894, S0=>nx36053);
   ix7895 : nor02ii port map ( Y=>nx7894, A0=>nx27299, A1=>nx36059);
   ix7889 : xor2 port map ( Y=>nx13153, A0=>nx27314, A1=>nx27545);
   ix27331 : or02 port map ( Y=>nx27330, A0=>nx27267, A1=>nx35761);
   ix7877 : xor2 port map ( Y=>nx13155, A0=>nx27348, A1=>nx35341);
   ix18494 : mux21_ni port map ( Y=>nx18493, A0=>
      booth_booth_integrtaion_9_booth_output_20, A1=>nx7870, S0=>nx36053);
   ix7871 : nor02ii port map ( Y=>nx7870, A0=>nx27336, A1=>nx36059);
   ix7865 : xor2 port map ( Y=>nx13157, A0=>nx27353, A1=>nx27542);
   ix7853 : xor2 port map ( Y=>nx13159, A0=>nx27383, A1=>nx35343);
   ix18474 : mux21_ni port map ( Y=>nx18473, A0=>
      booth_booth_integrtaion_9_booth_output_22, A1=>nx7846, S0=>nx36053);
   ix7847 : nor02ii port map ( Y=>nx7846, A0=>nx27371, A1=>nx36059);
   ix7841 : xor2 port map ( Y=>nx13161, A0=>nx27388, A1=>nx27539);
   ix7829 : xor2 port map ( Y=>nx13162, A0=>nx27418, A1=>nx35345);
   ix18454 : mux21_ni port map ( Y=>nx18453, A0=>
      booth_booth_integrtaion_9_booth_output_24, A1=>nx7822, S0=>nx36053);
   ix7823 : nor02ii port map ( Y=>nx7822, A0=>nx27406, A1=>nx36061);
   ix7817 : xor2 port map ( Y=>nx13163, A0=>nx27423, A1=>nx27536);
   ix7805 : xor2 port map ( Y=>nx13165, A0=>nx27453, A1=>nx35347);
   ix18434 : mux21_ni port map ( Y=>nx18433, A0=>
      booth_booth_integrtaion_9_booth_output_26, A1=>nx7798, S0=>nx36053);
   ix7799 : nor02ii port map ( Y=>nx7798, A0=>nx27441, A1=>nx36061);
   ix7793 : xor2 port map ( Y=>nx13167, A0=>nx27458, A1=>nx27533);
   ix7781 : xor2 port map ( Y=>nx13169, A0=>nx27488, A1=>nx35349);
   ix18414 : mux21_ni port map ( Y=>nx18413, A0=>
      booth_booth_integrtaion_9_booth_output_28, A1=>nx7774, S0=>nx35331);
   ix7775 : nor02ii port map ( Y=>nx7774, A0=>nx27476, A1=>nx36061);
   ix7769 : xor2 port map ( Y=>nx13170, A0=>nx27493, A1=>nx27530);
   ix7757 : xor2 port map ( Y=>nx13171, A0=>nx27523, A1=>nx35351);
   ix18394 : mux21_ni port map ( Y=>nx18393, A0=>
      booth_booth_integrtaion_9_booth_output_31, A1=>nx7750, S0=>nx35331);
   ix7751 : nor02ii port map ( Y=>nx7750, A0=>nx27511, A1=>nx36061);
   ix7745 : xor2 port map ( Y=>nx7744, A0=>nx27523, A1=>nx27526);
   ix7931 : nor02ii port map ( Y=>nx7930, A0=>nx7394, A1=>nx36061);
   ix27577 : or03 port map ( Y=>nx27576, A0=>nx27760, A1=>nx35843, A2=>
      nx35361);
   ix18984 : mux21_ni port map ( Y=>nx18983, A0=>label_10_output(14), A1=>
      label_10_input_14, S0=>nx36241);
   ix8575 : mux21_ni port map ( Y=>nx8574, A0=>nx8570, A1=>
      label_10_input_state_machine_14, S0=>nx35919);
   ix18164 : mux21_ni port map ( Y=>nx18163, A0=>
      label_10_input_state_machine_14, A1=>mdr_data_out(158), S0=>nx36201);
   ix18974 : mux21_ni port map ( Y=>nx18973, A0=>label_10_output(13), A1=>
      label_10_input_13, S0=>nx36241);
   ix8549 : mux21_ni port map ( Y=>nx8548, A0=>nx8544, A1=>
      label_10_input_state_machine_13, S0=>nx35921);
   ix18964 : mux21_ni port map ( Y=>nx18963, A0=>
      label_10_input_state_machine_13, A1=>mdr_data_out(157), S0=>nx36201);
   ix18934 : mux21_ni port map ( Y=>nx18933, A0=>label_10_output(11), A1=>
      label_10_input_11, S0=>nx36241);
   ix8485 : mux21_ni port map ( Y=>nx8484, A0=>nx8480, A1=>
      label_10_input_state_machine_11, S0=>nx35921);
   ix18924 : mux21_ni port map ( Y=>nx18923, A0=>
      label_10_input_state_machine_11, A1=>mdr_data_out(155), S0=>nx36203);
   ix18894 : mux21_ni port map ( Y=>nx18893, A0=>label_10_output(9), A1=>
      label_10_input_9, S0=>nx36241);
   ix8421 : mux21_ni port map ( Y=>nx8420, A0=>nx8416, A1=>
      label_10_input_state_machine_9, S0=>nx35921);
   ix18884 : mux21_ni port map ( Y=>nx18883, A0=>
      label_10_input_state_machine_9, A1=>mdr_data_out(153), S0=>nx36203);
   ix18854 : mux21_ni port map ( Y=>nx18853, A0=>label_10_output(7), A1=>
      label_10_input_7, S0=>nx36243);
   ix8357 : mux21_ni port map ( Y=>nx8356, A0=>nx8352, A1=>
      label_10_input_state_machine_7, S0=>nx35921);
   ix18844 : mux21_ni port map ( Y=>nx18843, A0=>
      label_10_input_state_machine_7, A1=>mdr_data_out(151), S0=>nx36203);
   ix18814 : mux21_ni port map ( Y=>nx18813, A0=>label_10_output(5), A1=>
      label_10_input_5, S0=>nx36243);
   ix8293 : mux21_ni port map ( Y=>nx8292, A0=>nx8288, A1=>
      label_10_input_state_machine_5, S0=>nx35921);
   ix18804 : mux21_ni port map ( Y=>nx18803, A0=>
      label_10_input_state_machine_5, A1=>mdr_data_out(149), S0=>nx36203);
   ix18774 : mux21_ni port map ( Y=>nx18773, A0=>label_10_output(3), A1=>
      label_10_input_3, S0=>nx36243);
   ix8229 : mux21_ni port map ( Y=>nx8228, A0=>nx8224, A1=>
      label_10_input_state_machine_3, S0=>nx35921);
   ix18764 : mux21_ni port map ( Y=>nx18763, A0=>
      label_10_input_state_machine_3, A1=>mdr_data_out(147), S0=>nx36203);
   ix18734 : mux21_ni port map ( Y=>nx18733, A0=>label_10_output(1), A1=>
      label_10_input_1, S0=>nx36243);
   ix8165 : mux21_ni port map ( Y=>nx8164, A0=>nx8160, A1=>
      label_10_input_state_machine_1, S0=>nx35921);
   ix18724 : mux21_ni port map ( Y=>nx18723, A0=>
      label_10_input_state_machine_1, A1=>mdr_data_out(145), S0=>nx36203);
   ix27669 : xnor2 port map ( Y=>nx27668, A0=>nx27566, A1=>nx27678);
   ix18754 : mux21_ni port map ( Y=>nx18753, A0=>label_10_output(2), A1=>
      label_10_input_2, S0=>nx36243);
   ix8197 : mux21_ni port map ( Y=>nx8196, A0=>nx8192, A1=>
      label_10_input_state_machine_2, S0=>nx35923);
   ix18744 : mux21_ni port map ( Y=>nx18743, A0=>
      label_10_input_state_machine_2, A1=>mdr_data_out(146), S0=>nx36203);
   ix27684 : xnor2 port map ( Y=>nx27683, A0=>nx27564, A1=>nx27693);
   ix18794 : mux21_ni port map ( Y=>nx18793, A0=>label_10_output(4), A1=>
      label_10_input_4, S0=>nx36243);
   ix8261 : mux21_ni port map ( Y=>nx8260, A0=>nx8256, A1=>
      label_10_input_state_machine_4, S0=>nx35923);
   ix18784 : mux21_ni port map ( Y=>nx18783, A0=>
      label_10_input_state_machine_4, A1=>mdr_data_out(148), S0=>nx36205);
   ix27699 : xnor2 port map ( Y=>nx27698, A0=>nx27562, A1=>nx27708);
   ix18834 : mux21_ni port map ( Y=>nx18833, A0=>label_10_output(6), A1=>
      label_10_input_6, S0=>nx36243);
   ix8325 : mux21_ni port map ( Y=>nx8324, A0=>nx8320, A1=>
      label_10_input_state_machine_6, S0=>nx35923);
   ix18824 : mux21_ni port map ( Y=>nx18823, A0=>
      label_10_input_state_machine_6, A1=>mdr_data_out(150), S0=>nx36205);
   ix27714 : xnor2 port map ( Y=>nx27713, A0=>nx27560, A1=>nx27723);
   ix18874 : mux21_ni port map ( Y=>nx18873, A0=>label_10_output(8), A1=>
      label_10_input_8, S0=>nx36245);
   ix8389 : mux21_ni port map ( Y=>nx8388, A0=>nx8384, A1=>
      label_10_input_state_machine_8, S0=>nx35923);
   ix18864 : mux21_ni port map ( Y=>nx18863, A0=>
      label_10_input_state_machine_8, A1=>mdr_data_out(152), S0=>nx36205);
   ix27729 : xnor2 port map ( Y=>nx27728, A0=>nx27558, A1=>nx27738);
   ix18914 : mux21_ni port map ( Y=>nx18913, A0=>label_10_output(10), A1=>
      label_10_input_10, S0=>nx36245);
   ix8453 : mux21_ni port map ( Y=>nx8452, A0=>nx8448, A1=>
      label_10_input_state_machine_10, S0=>nx35923);
   ix18904 : mux21_ni port map ( Y=>nx18903, A0=>
      label_10_input_state_machine_10, A1=>mdr_data_out(154), S0=>nx36205);
   ix27744 : xnor2 port map ( Y=>nx27743, A0=>nx27556, A1=>nx27753);
   ix18954 : mux21_ni port map ( Y=>nx18953, A0=>label_10_output(12), A1=>
      label_10_input_12, S0=>nx36245);
   ix8517 : mux21_ni port map ( Y=>nx8516, A0=>nx8512, A1=>
      label_10_input_state_machine_12, S0=>nx35923);
   ix18944 : mux21_ni port map ( Y=>nx18943, A0=>
      label_10_input_state_machine_12, A1=>mdr_data_out(156), S0=>nx36205);
   ix27759 : xnor2 port map ( Y=>nx27758, A0=>nx27554, A1=>nx27760);
   ix27766 : or03 port map ( Y=>nx27765, A0=>nx27949, A1=>nx35843, A2=>
      nx35361);
   ix19274 : mux21_ni port map ( Y=>nx19273, A0=>label_9_output(14), A1=>
      label_9_input_14, S0=>nx36245);
   ix9025 : mux21_ni port map ( Y=>nx9024, A0=>nx9020, A1=>
      label_9_input_state_machine_14, S0=>nx35925);
   ix19004 : mux21_ni port map ( Y=>nx19003, A0=>
      label_9_input_state_machine_14, A1=>mdr_data_out(142), S0=>nx36205);
   ix19264 : mux21_ni port map ( Y=>nx19263, A0=>label_9_output(13), A1=>
      label_9_input_13, S0=>nx36245);
   ix8999 : mux21_ni port map ( Y=>nx8998, A0=>nx8994, A1=>
      label_9_input_state_machine_13, S0=>nx35925);
   ix19254 : mux21_ni port map ( Y=>nx19253, A0=>
      label_9_input_state_machine_13, A1=>mdr_data_out(141), S0=>nx36205);
   ix19224 : mux21_ni port map ( Y=>nx19223, A0=>label_9_output(11), A1=>
      label_9_input_11, S0=>nx36245);
   ix8935 : mux21_ni port map ( Y=>nx8934, A0=>nx8930, A1=>
      label_9_input_state_machine_11, S0=>nx35925);
   ix19214 : mux21_ni port map ( Y=>nx19213, A0=>
      label_9_input_state_machine_11, A1=>mdr_data_out(139), S0=>nx36207);
   ix19184 : mux21_ni port map ( Y=>nx19183, A0=>label_9_output(9), A1=>
      label_9_input_9, S0=>nx36245);
   ix8871 : mux21_ni port map ( Y=>nx8870, A0=>nx8866, A1=>
      label_9_input_state_machine_9, S0=>nx35925);
   ix19174 : mux21_ni port map ( Y=>nx19173, A0=>
      label_9_input_state_machine_9, A1=>mdr_data_out(137), S0=>nx36207);
   ix19144 : mux21_ni port map ( Y=>nx19143, A0=>label_9_output(7), A1=>
      label_9_input_7, S0=>nx36247);
   ix8807 : mux21_ni port map ( Y=>nx8806, A0=>nx8802, A1=>
      label_9_input_state_machine_7, S0=>nx35923);
   ix19134 : mux21_ni port map ( Y=>nx19133, A0=>
      label_9_input_state_machine_7, A1=>mdr_data_out(135), S0=>nx36207);
   ix19104 : mux21_ni port map ( Y=>nx19103, A0=>label_9_output(5), A1=>
      label_9_input_5, S0=>nx36247);
   ix8743 : mux21_ni port map ( Y=>nx8742, A0=>nx8738, A1=>
      label_9_input_state_machine_5, S0=>nx35165);
   ix19094 : mux21_ni port map ( Y=>nx19093, A0=>
      label_9_input_state_machine_5, A1=>mdr_data_out(133), S0=>nx36207);
   ix19064 : mux21_ni port map ( Y=>nx19063, A0=>label_9_output(3), A1=>
      label_9_input_3, S0=>nx36247);
   ix8679 : mux21_ni port map ( Y=>nx8678, A0=>nx8674, A1=>
      label_9_input_state_machine_3, S0=>nx35165);
   ix19054 : mux21_ni port map ( Y=>nx19053, A0=>
      label_9_input_state_machine_3, A1=>mdr_data_out(131), S0=>nx36207);
   ix19024 : mux21_ni port map ( Y=>nx19023, A0=>label_9_output(1), A1=>
      label_9_input_1, S0=>nx36247);
   ix8615 : mux21_ni port map ( Y=>nx8614, A0=>nx8610, A1=>
      label_9_input_state_machine_1, S0=>nx35165);
   ix19014 : mux21_ni port map ( Y=>nx19013, A0=>
      label_9_input_state_machine_1, A1=>mdr_data_out(129), S0=>nx36207);
   ix27858 : xnor2 port map ( Y=>nx27857, A0=>nx27127, A1=>nx27867);
   ix19044 : mux21_ni port map ( Y=>nx19043, A0=>label_9_output(2), A1=>
      label_9_input_2, S0=>nx36247);
   ix8647 : mux21_ni port map ( Y=>nx8646, A0=>nx8642, A1=>
      label_9_input_state_machine_2, S0=>nx35165);
   ix19034 : mux21_ni port map ( Y=>nx19033, A0=>
      label_9_input_state_machine_2, A1=>mdr_data_out(130), S0=>nx36207);
   ix27873 : xnor2 port map ( Y=>nx27872, A0=>nx27125, A1=>nx27882);
   ix19084 : mux21_ni port map ( Y=>nx19083, A0=>label_9_output(4), A1=>
      label_9_input_4, S0=>nx36247);
   ix8711 : mux21_ni port map ( Y=>nx8710, A0=>nx8706, A1=>
      label_9_input_state_machine_4, S0=>nx35165);
   ix19074 : mux21_ni port map ( Y=>nx19073, A0=>
      label_9_input_state_machine_4, A1=>mdr_data_out(132), S0=>nx36209);
   ix27888 : xnor2 port map ( Y=>nx27887, A0=>nx27123, A1=>nx27897);
   ix19124 : mux21_ni port map ( Y=>nx19123, A0=>label_9_output(6), A1=>
      label_9_input_6, S0=>nx36247);
   ix8775 : mux21_ni port map ( Y=>nx8774, A0=>nx8770, A1=>
      label_9_input_state_machine_6, S0=>nx35165);
   ix19114 : mux21_ni port map ( Y=>nx19113, A0=>
      label_9_input_state_machine_6, A1=>mdr_data_out(134), S0=>nx36209);
   ix27903 : xnor2 port map ( Y=>nx27902, A0=>nx27121, A1=>nx27912);
   ix19164 : mux21_ni port map ( Y=>nx19163, A0=>label_9_output(8), A1=>
      label_9_input_8, S0=>nx36249);
   ix8839 : mux21_ni port map ( Y=>nx8838, A0=>nx8834, A1=>
      label_9_input_state_machine_8, S0=>nx35165);
   ix19154 : mux21_ni port map ( Y=>nx19153, A0=>
      label_9_input_state_machine_8, A1=>mdr_data_out(136), S0=>nx36209);
   ix27918 : xnor2 port map ( Y=>nx27917, A0=>nx27119, A1=>nx27927);
   ix19204 : mux21_ni port map ( Y=>nx19203, A0=>label_9_output(10), A1=>
      label_9_input_10, S0=>nx36249);
   ix8903 : mux21_ni port map ( Y=>nx8902, A0=>nx8898, A1=>
      label_9_input_state_machine_10, S0=>nx35925);
   ix19194 : mux21_ni port map ( Y=>nx19193, A0=>
      label_9_input_state_machine_10, A1=>mdr_data_out(138), S0=>nx36209);
   ix27933 : xnor2 port map ( Y=>nx27932, A0=>nx27117, A1=>nx27942);
   ix19244 : mux21_ni port map ( Y=>nx19243, A0=>label_9_output(12), A1=>
      label_9_input_12, S0=>nx36249);
   ix8967 : mux21_ni port map ( Y=>nx8966, A0=>nx8962, A1=>
      label_9_input_state_machine_12, S0=>nx35927);
   ix19234 : mux21_ni port map ( Y=>nx19233, A0=>
      label_9_input_state_machine_12, A1=>mdr_data_out(140), S0=>nx36209);
   ix27948 : xnor2 port map ( Y=>nx27947, A0=>nx27115, A1=>nx27949);
   ix9045 : xnor2 port map ( Y=>nx9044, A0=>nx27573, A1=>nx27763);
   ix27953 : xnor2 port map ( Y=>nx27952, A0=>nx27956, A1=>
      max_calc_comparator_fifth_inp1_13);
   ix27971 : or03 port map ( Y=>nx27970, A0=>nx27753, A1=>nx35845, A2=>
      nx35361);
   ix27977 : or03 port map ( Y=>nx27976, A0=>nx27942, A1=>nx35845, A2=>
      nx35361);
   ix9081 : xnor2 port map ( Y=>nx9080, A0=>nx27967, A1=>nx27974);
   ix27981 : xnor2 port map ( Y=>nx27980, A0=>nx27984, A1=>
      max_calc_comparator_fifth_inp1_11);
   ix27999 : or03 port map ( Y=>nx27998, A0=>nx27738, A1=>nx35845, A2=>
      nx36065);
   ix28005 : or03 port map ( Y=>nx28004, A0=>nx27927, A1=>nx35845, A2=>
      nx36065);
   ix9117 : xnor2 port map ( Y=>nx9116, A0=>nx27995, A1=>nx28002);
   ix28009 : xnor2 port map ( Y=>nx28008, A0=>nx28012, A1=>
      max_calc_comparator_fifth_inp1_9);
   ix28027 : or03 port map ( Y=>nx28026, A0=>nx27723, A1=>nx35845, A2=>
      nx36065);
   ix28033 : or03 port map ( Y=>nx28032, A0=>nx27912, A1=>nx35845, A2=>
      nx36065);
   ix9153 : xnor2 port map ( Y=>nx9152, A0=>nx28023, A1=>nx28030);
   ix28037 : xnor2 port map ( Y=>nx28036, A0=>nx28040, A1=>
      max_calc_comparator_fifth_inp1_7);
   ix28055 : or03 port map ( Y=>nx28054, A0=>nx27708, A1=>nx35845, A2=>
      nx36065);
   ix28061 : or03 port map ( Y=>nx28060, A0=>nx27897, A1=>nx35847, A2=>
      nx36065);
   ix9189 : xnor2 port map ( Y=>nx9188, A0=>nx28051, A1=>nx28058);
   ix28065 : xnor2 port map ( Y=>nx28064, A0=>nx28068, A1=>
      max_calc_comparator_fifth_inp1_5);
   ix28083 : or03 port map ( Y=>nx28082, A0=>nx27693, A1=>nx35847, A2=>
      nx36065);
   ix28089 : or03 port map ( Y=>nx28088, A0=>nx27882, A1=>nx35847, A2=>
      nx35363);
   ix9225 : xnor2 port map ( Y=>nx9224, A0=>nx28079, A1=>nx28086);
   ix28093 : xnor2 port map ( Y=>nx28092, A0=>nx28096, A1=>
      max_calc_comparator_fifth_inp1_3);
   ix28111 : or03 port map ( Y=>nx28110, A0=>nx27678, A1=>nx35847, A2=>
      nx35363);
   ix28117 : or03 port map ( Y=>nx28116, A0=>nx27867, A1=>nx35847, A2=>
      nx35363);
   ix9261 : xnor2 port map ( Y=>nx9260, A0=>nx28107, A1=>nx28114);
   ix9279 : xnor2 port map ( Y=>nx9278, A0=>nx28122, A1=>nx28126);
   ix9489 : xnor2 port map ( Y=>nx9488, A0=>nx28137, A1=>nx28155);
   ix19574 : mux21_ni port map ( Y=>nx19573, A0=>label_10_output(15), A1=>
      label_10_input_15, S0=>nx36249);
   ix9429 : mux21_ni port map ( Y=>nx9428, A0=>nx9424, A1=>
      label_10_input_state_machine_15, S0=>nx35927);
   ix19564 : mux21_ni port map ( Y=>nx19563, A0=>
      label_10_input_state_machine_15, A1=>mdr_data_out(159), S0=>nx36209);
   ix28151 : xor2 port map ( Y=>nx28150, A0=>nx27552, A1=>
      label_10_output(15));
   ix19604 : mux21_ni port map ( Y=>nx19603, A0=>label_9_output(15), A1=>
      label_9_input_15, S0=>nx36249);
   ix9469 : mux21_ni port map ( Y=>nx9468, A0=>nx9464, A1=>
      label_9_input_state_machine_15, S0=>nx35927);
   ix19594 : mux21_ni port map ( Y=>nx19593, A0=>
      label_9_input_state_machine_15, A1=>mdr_data_out(143), S0=>nx36209);
   ix28169 : xor2 port map ( Y=>nx28168, A0=>nx27113, A1=>label_9_output(15)
   );
   ix28173 : or04 port map ( Y=>nx28172, A0=>rst, A1=>nx26180, A2=>
      max_calc_state_3, A3=>nx26188);
   ix25474 : mux21_ni port map ( Y=>nx25473, A0=>
      max_calc_comparator_first_inp2_0, A1=>nx18892, S0=>nx36281);
   ix18893 : mux21_ni port map ( Y=>nx18892, A0=>nx18888, A1=>nx18864, S0=>
      nx35965);
   ix18865 : mux21_ni port map ( Y=>nx18864, A0=>max_calc_ans2_0, A1=>
      label_2_output(0), S0=>nx35987);
   ix16374 : mux21_ni port map ( Y=>nx16373, A0=>label_2_output(0), A1=>
      label_2_input_0, S0=>nx36249);
   ix16364 : mux21_ni port map ( Y=>nx16363, A0=>
      label_2_input_state_machine_0, A1=>mdr_data_out(16), S0=>nx36211);
   ix16354 : mux21_ni port map ( Y=>nx16353, A0=>nx35727, A1=>nx4398, S0=>
      nx35379);
   ix4399 : mux21_ni port map ( Y=>nx4398, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_1_1, S0=>nx36085);
   ix16344 : mux21_ni port map ( Y=>nx16343, A0=>
      booth_booth_integration_output_1_1, A1=>nx4386, S0=>nx35379);
   ix4387 : mux21_ni port map ( Y=>nx4386, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_1_2, S0=>nx36085);
   ix16334 : mux21_ni port map ( Y=>nx16333, A0=>
      booth_booth_integration_output_1_2, A1=>nx4374, S0=>nx35379);
   ix4375 : mux21_ni port map ( Y=>nx4374, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_1_3, S0=>nx36085);
   ix16324 : mux21_ni port map ( Y=>nx16323, A0=>
      booth_booth_integration_output_1_3, A1=>nx4362, S0=>nx35379);
   ix4363 : mux21_ni port map ( Y=>nx4362, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_1_4, S0=>nx36085);
   ix16314 : mux21_ni port map ( Y=>nx16313, A0=>
      booth_booth_integration_output_1_4, A1=>nx4350, S0=>nx35379);
   ix4351 : mux21_ni port map ( Y=>nx4350, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_1_5, S0=>nx36085);
   ix16304 : mux21_ni port map ( Y=>nx16303, A0=>
      booth_booth_integration_output_1_5, A1=>nx4338, S0=>nx35379);
   ix4339 : mux21_ni port map ( Y=>nx4338, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_1_6, S0=>nx36087);
   ix16294 : mux21_ni port map ( Y=>nx16293, A0=>
      booth_booth_integration_output_1_6, A1=>nx4326, S0=>nx35379);
   ix4327 : mux21_ni port map ( Y=>nx4326, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_1_7, S0=>nx36087);
   ix16284 : mux21_ni port map ( Y=>nx16283, A0=>
      booth_booth_integration_output_1_7, A1=>nx4314, S0=>nx36077);
   ix4315 : mux21_ni port map ( Y=>nx4314, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_1_8, S0=>nx36087);
   ix16274 : mux21_ni port map ( Y=>nx16273, A0=>
      booth_booth_integration_output_1_8, A1=>nx4302, S0=>nx36077);
   ix4303 : mux21_ni port map ( Y=>nx4302, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_1_9, S0=>nx36087);
   ix16264 : mux21_ni port map ( Y=>nx16263, A0=>
      booth_booth_integration_output_1_9, A1=>nx4290, S0=>nx36077);
   ix4291 : mux21_ni port map ( Y=>nx4290, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_1_10, S0=>nx36087);
   ix16254 : mux21_ni port map ( Y=>nx16253, A0=>
      booth_booth_integration_output_1_10, A1=>nx4278, S0=>nx36079);
   ix4279 : mux21_ni port map ( Y=>nx4278, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_1_11, S0=>nx36087);
   ix16244 : mux21_ni port map ( Y=>nx16243, A0=>
      booth_booth_integration_output_1_11, A1=>nx4266, S0=>nx36079);
   ix4267 : mux21_ni port map ( Y=>nx4266, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_1_12, S0=>nx36087);
   ix16234 : mux21_ni port map ( Y=>nx16233, A0=>
      booth_booth_integration_output_1_12, A1=>nx4254, S0=>nx36079);
   ix4255 : mux21_ni port map ( Y=>nx4254, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_1_13, S0=>nx36089);
   ix16224 : mux21_ni port map ( Y=>nx16223, A0=>
      booth_booth_integration_output_1_13, A1=>nx4242, S0=>nx36079);
   ix4243 : mux21_ni port map ( Y=>nx4242, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_1_14, S0=>nx36089);
   ix16214 : mux21_ni port map ( Y=>nx16213, A0=>
      booth_booth_integration_output_1_14, A1=>nx4230, S0=>nx36079);
   ix4231 : mux21_ni port map ( Y=>nx4230, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_1_15, S0=>nx36089);
   ix16204 : mux21 port map ( Y=>nx16203, A0=>nx28594, A1=>nx28236, S0=>
      nx36079);
   ix15854 : mux21_ni port map ( Y=>nx15853, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_0, A1=>nx34635, S0=>nx35815
   );
   ix15840 : and02 port map ( Y=>nx15839, A0=>nx36323, A1=>
      booth_booth_integrtaion_1_shift_Reg_count_0);
   ix16034 : mux21_ni port map ( Y=>nx16033, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_9, A1=>nx34621, S0=>nx35815
   );
   ix16024 : mux21_ni port map ( Y=>nx16023, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_8, S0=>nx36079);
   ix16014 : mux21_ni port map ( Y=>nx16013, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_8, S0=>nx35815);
   ix16004 : mux21_ni port map ( Y=>nx16003, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_7, S0=>nx36081);
   ix15994 : mux21_ni port map ( Y=>nx15993, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_7, S0=>nx35815);
   ix15984 : mux21_ni port map ( Y=>nx15983, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_6, S0=>nx36081);
   ix15974 : mux21_ni port map ( Y=>nx15973, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_6, S0=>nx35815);
   ix15964 : mux21_ni port map ( Y=>nx15963, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_5, S0=>nx36081);
   ix15954 : mux21_ni port map ( Y=>nx15953, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_5, S0=>nx35815);
   ix15944 : mux21_ni port map ( Y=>nx15943, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_4, S0=>nx36081);
   ix15934 : mux21_ni port map ( Y=>nx15933, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_4, S0=>nx35817);
   ix15924 : mux21_ni port map ( Y=>nx15923, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_3, S0=>nx36081);
   ix15914 : mux21_ni port map ( Y=>nx15913, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_3, S0=>nx35817);
   ix15904 : mux21_ni port map ( Y=>nx15903, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_2, S0=>nx36081);
   ix15894 : mux21_ni port map ( Y=>nx15893, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_2, S0=>nx35817);
   ix15884 : mux21_ni port map ( Y=>nx15883, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_1, S0=>nx36081);
   ix15874 : mux21_ni port map ( Y=>nx15873, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_1_shift_Reg_output_1, S0=>nx35817);
   ix15864 : mux21_ni port map ( Y=>nx15863, A0=>
      booth_booth_integrtaion_1_shift_Reg_count_1, A1=>nx34635, S0=>nx36083
   );
   ix3671 : and02 port map ( Y=>nx3670, A0=>nx28309, A1=>nx35727);
   ix28312 : or03 port map ( Y=>nx28311, A0=>nx28313, A1=>
      booth_booth_integrtaion_1_shift_reg_output_0, A2=>nx36323);
   ix16194 : mux21_ni port map ( Y=>nx16193, A0=>
      booth_booth_integrtaion_1_booth_output_16, A1=>nx4200, S0=>nx36083);
   ix4201 : nor02ii port map ( Y=>nx4200, A0=>nx28320, A1=>nx36089);
   ix3677 : nor02ii port map ( Y=>nx3676, A0=>nx28304, A1=>
      booth_booth_integrtaion_1_booth_output_16);
   ix4195 : xor2 port map ( Y=>nx13017, A0=>nx28326, A1=>nx28590);
   ix4183 : xor2 port map ( Y=>nx13018, A0=>nx28351, A1=>nx35385);
   ix16174 : mux21_ni port map ( Y=>nx16173, A0=>
      booth_booth_integrtaion_1_booth_output_18, A1=>nx4176, S0=>nx36083);
   ix4177 : nor02ii port map ( Y=>nx4176, A0=>nx28341, A1=>nx36089);
   ix4171 : xor2 port map ( Y=>nx13019, A0=>nx28356, A1=>nx28587);
   ix28373 : or02 port map ( Y=>nx28372, A0=>nx28309, A1=>nx35729);
   ix4159 : xor2 port map ( Y=>nx13021, A0=>nx28390, A1=>nx35387);
   ix16154 : mux21_ni port map ( Y=>nx16153, A0=>
      booth_booth_integrtaion_1_booth_output_20, A1=>nx4152, S0=>nx36083);
   ix4153 : nor02ii port map ( Y=>nx4152, A0=>nx28378, A1=>nx36089);
   ix4147 : xor2 port map ( Y=>nx13023, A0=>nx28395, A1=>nx28584);
   ix4135 : xor2 port map ( Y=>nx13025, A0=>nx28425, A1=>nx35389);
   ix16134 : mux21_ni port map ( Y=>nx16133, A0=>
      booth_booth_integrtaion_1_booth_output_22, A1=>nx4128, S0=>nx36083);
   ix4129 : nor02ii port map ( Y=>nx4128, A0=>nx28413, A1=>nx36089);
   ix4123 : xor2 port map ( Y=>nx13026, A0=>nx28430, A1=>nx28581);
   ix4111 : xor2 port map ( Y=>nx13027, A0=>nx28460, A1=>nx35391);
   ix16114 : mux21_ni port map ( Y=>nx16113, A0=>
      booth_booth_integrtaion_1_booth_output_24, A1=>nx4104, S0=>nx36083);
   ix4105 : nor02ii port map ( Y=>nx4104, A0=>nx28448, A1=>nx36091);
   ix4099 : xor2 port map ( Y=>nx13029, A0=>nx28465, A1=>nx28578);
   ix4087 : xor2 port map ( Y=>nx13031, A0=>nx28495, A1=>nx35393);
   ix16094 : mux21_ni port map ( Y=>nx16093, A0=>
      booth_booth_integrtaion_1_booth_output_26, A1=>nx4080, S0=>nx36083);
   ix4081 : nor02ii port map ( Y=>nx4080, A0=>nx28483, A1=>nx36091);
   ix4075 : xor2 port map ( Y=>nx13033, A0=>nx28500, A1=>nx28575);
   ix4063 : xor2 port map ( Y=>nx13035, A0=>nx28530, A1=>nx35395);
   ix16074 : mux21_ni port map ( Y=>nx16073, A0=>
      booth_booth_integrtaion_1_booth_output_28, A1=>nx4056, S0=>nx35377);
   ix4057 : nor02ii port map ( Y=>nx4056, A0=>nx28518, A1=>nx36091);
   ix4051 : xor2 port map ( Y=>nx13037, A0=>nx28535, A1=>nx28572);
   ix4039 : xor2 port map ( Y=>nx13039, A0=>nx28565, A1=>nx35397);
   ix16054 : mux21_ni port map ( Y=>nx16053, A0=>
      booth_booth_integrtaion_1_booth_output_31, A1=>nx4032, S0=>nx35377);
   ix4033 : nor02ii port map ( Y=>nx4032, A0=>nx28553, A1=>nx36091);
   ix4027 : xor2 port map ( Y=>nx4026, A0=>nx28565, A1=>nx28568);
   ix4213 : nor02ii port map ( Y=>nx4212, A0=>nx3676, A1=>nx36091);
   ix25444 : mux21_ni port map ( Y=>nx25443, A0=>nx18854, A1=>
      max_calc_ans2_0, S0=>nx35851);
   ix18855 : mux21 port map ( Y=>nx18854, A0=>nx30546, A1=>nx28617, S0=>
      nx35899);
   ix16933 : mux21_ni port map ( Y=>nx16932, A0=>max_calc_ans3_0, A1=>
      label_3_output(0), S0=>nx35977);
   ix15524 : mux21_ni port map ( Y=>nx15523, A0=>label_3_output(0), A1=>
      label_3_input_0, S0=>nx36249);
   ix15514 : mux21_ni port map ( Y=>nx15513, A0=>
      label_3_input_state_machine_0, A1=>mdr_data_out(32), S0=>nx36211);
   ix15504 : mux21_ni port map ( Y=>nx15503, A0=>nx35723, A1=>nx3060, S0=>
      nx35405);
   ix3061 : mux21_ni port map ( Y=>nx3060, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_2_1, S0=>nx36101);
   ix15494 : mux21_ni port map ( Y=>nx15493, A0=>
      booth_booth_integration_output_2_1, A1=>nx3048, S0=>nx35405);
   ix3049 : mux21_ni port map ( Y=>nx3048, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_2_2, S0=>nx36101);
   ix15484 : mux21_ni port map ( Y=>nx15483, A0=>
      booth_booth_integration_output_2_2, A1=>nx3036, S0=>nx35405);
   ix3037 : mux21_ni port map ( Y=>nx3036, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_2_3, S0=>nx36101);
   ix15474 : mux21_ni port map ( Y=>nx15473, A0=>
      booth_booth_integration_output_2_3, A1=>nx3024, S0=>nx35405);
   ix3025 : mux21_ni port map ( Y=>nx3024, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_2_4, S0=>nx36101);
   ix15464 : mux21_ni port map ( Y=>nx15463, A0=>
      booth_booth_integration_output_2_4, A1=>nx3012, S0=>nx35405);
   ix3013 : mux21_ni port map ( Y=>nx3012, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_2_5, S0=>nx36101);
   ix15454 : mux21_ni port map ( Y=>nx15453, A0=>
      booth_booth_integration_output_2_5, A1=>nx3000, S0=>nx35405);
   ix3001 : mux21_ni port map ( Y=>nx3000, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_2_6, S0=>nx36103);
   ix15444 : mux21_ni port map ( Y=>nx15443, A0=>
      booth_booth_integration_output_2_6, A1=>nx2988, S0=>nx35405);
   ix2989 : mux21_ni port map ( Y=>nx2988, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_2_7, S0=>nx36103);
   ix15434 : mux21_ni port map ( Y=>nx15433, A0=>
      booth_booth_integration_output_2_7, A1=>nx2976, S0=>nx36093);
   ix2977 : mux21_ni port map ( Y=>nx2976, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_2_8, S0=>nx36103);
   ix15424 : mux21_ni port map ( Y=>nx15423, A0=>
      booth_booth_integration_output_2_8, A1=>nx2964, S0=>nx36093);
   ix2965 : mux21_ni port map ( Y=>nx2964, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_2_9, S0=>nx36103);
   ix15414 : mux21_ni port map ( Y=>nx15413, A0=>
      booth_booth_integration_output_2_9, A1=>nx2952, S0=>nx36093);
   ix2953 : mux21_ni port map ( Y=>nx2952, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_2_10, S0=>nx36103);
   ix15404 : mux21_ni port map ( Y=>nx15403, A0=>
      booth_booth_integration_output_2_10, A1=>nx2940, S0=>nx36095);
   ix2941 : mux21_ni port map ( Y=>nx2940, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_2_11, S0=>nx36103);
   ix15394 : mux21_ni port map ( Y=>nx15393, A0=>
      booth_booth_integration_output_2_11, A1=>nx2928, S0=>nx36095);
   ix2929 : mux21_ni port map ( Y=>nx2928, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_2_12, S0=>nx36103);
   ix15384 : mux21_ni port map ( Y=>nx15383, A0=>
      booth_booth_integration_output_2_12, A1=>nx2916, S0=>nx36095);
   ix2917 : mux21_ni port map ( Y=>nx2916, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_2_13, S0=>nx36105);
   ix15374 : mux21_ni port map ( Y=>nx15373, A0=>
      booth_booth_integration_output_2_13, A1=>nx2904, S0=>nx36095);
   ix2905 : mux21_ni port map ( Y=>nx2904, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_2_14, S0=>nx36105);
   ix15364 : mux21_ni port map ( Y=>nx15363, A0=>
      booth_booth_integration_output_2_14, A1=>nx2892, S0=>nx36095);
   ix2893 : mux21_ni port map ( Y=>nx2892, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_2_15, S0=>nx36105);
   ix15354 : mux21 port map ( Y=>nx15353, A0=>nx29037, A1=>nx28679, S0=>
      nx36095);
   ix15004 : mux21_ni port map ( Y=>nx15003, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_0, A1=>nx34603, S0=>nx35819
   );
   ix14990 : and02 port map ( Y=>nx14989, A0=>nx36319, A1=>
      booth_booth_integrtaion_2_shift_Reg_count_0);
   ix15184 : mux21_ni port map ( Y=>nx15183, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_9, A1=>nx34589, S0=>nx35819
   );
   ix15174 : mux21_ni port map ( Y=>nx15173, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_8, S0=>nx36095);
   ix15164 : mux21_ni port map ( Y=>nx15163, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_8, S0=>nx35819);
   ix15154 : mux21_ni port map ( Y=>nx15153, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_7, S0=>nx36097);
   ix15144 : mux21_ni port map ( Y=>nx15143, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_7, S0=>nx35819);
   ix15134 : mux21_ni port map ( Y=>nx15133, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_6, S0=>nx36097);
   ix15124 : mux21_ni port map ( Y=>nx15123, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_6, S0=>nx35819);
   ix15114 : mux21_ni port map ( Y=>nx15113, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_5, S0=>nx36097);
   ix15104 : mux21_ni port map ( Y=>nx15103, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_5, S0=>nx35819);
   ix15094 : mux21_ni port map ( Y=>nx15093, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_4, S0=>nx36097);
   ix15084 : mux21_ni port map ( Y=>nx15083, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_4, S0=>nx35821);
   ix15074 : mux21_ni port map ( Y=>nx15073, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_3, S0=>nx36097);
   ix15064 : mux21_ni port map ( Y=>nx15063, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_3, S0=>nx35821);
   ix15054 : mux21_ni port map ( Y=>nx15053, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_2, S0=>nx36097);
   ix15044 : mux21_ni port map ( Y=>nx15043, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_2, S0=>nx35821);
   ix15034 : mux21_ni port map ( Y=>nx15033, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_1, S0=>nx36097);
   ix15024 : mux21_ni port map ( Y=>nx15023, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_2_shift_Reg_output_1, S0=>nx35821);
   ix15014 : mux21_ni port map ( Y=>nx15013, A0=>
      booth_booth_integrtaion_2_shift_Reg_count_1, A1=>nx34603, S0=>nx36099
   );
   ix2333 : and02 port map ( Y=>nx2332, A0=>nx28752, A1=>nx35723);
   ix28755 : or03 port map ( Y=>nx28754, A0=>nx28756, A1=>
      booth_booth_integrtaion_2_shift_reg_output_0, A2=>nx36319);
   ix15344 : mux21_ni port map ( Y=>nx15343, A0=>
      booth_booth_integrtaion_2_booth_output_16, A1=>nx2862, S0=>nx36099);
   ix2863 : nor02ii port map ( Y=>nx2862, A0=>nx28763, A1=>nx36105);
   ix2339 : nor02ii port map ( Y=>nx2338, A0=>nx28747, A1=>
      booth_booth_integrtaion_2_booth_output_16);
   ix2857 : xor2 port map ( Y=>nx12965, A0=>nx28769, A1=>nx29033);
   ix2845 : xor2 port map ( Y=>nx12967, A0=>nx28794, A1=>nx35411);
   ix15324 : mux21_ni port map ( Y=>nx15323, A0=>
      booth_booth_integrtaion_2_booth_output_18, A1=>nx2838, S0=>nx36099);
   ix2839 : nor02ii port map ( Y=>nx2838, A0=>nx28784, A1=>nx36105);
   ix2833 : xor2 port map ( Y=>nx12969, A0=>nx28799, A1=>nx29030);
   ix28816 : or02 port map ( Y=>nx28815, A0=>nx28752, A1=>nx35725);
   ix2821 : xor2 port map ( Y=>nx12970, A0=>nx28833, A1=>nx35413);
   ix15304 : mux21_ni port map ( Y=>nx15303, A0=>
      booth_booth_integrtaion_2_booth_output_20, A1=>nx2814, S0=>nx36099);
   ix2815 : nor02ii port map ( Y=>nx2814, A0=>nx28821, A1=>nx36105);
   ix2809 : xor2 port map ( Y=>nx12971, A0=>nx28838, A1=>nx29027);
   ix2797 : xor2 port map ( Y=>nx12973, A0=>nx28868, A1=>nx35415);
   ix15284 : mux21_ni port map ( Y=>nx15283, A0=>
      booth_booth_integrtaion_2_booth_output_22, A1=>nx2790, S0=>nx36099);
   ix2791 : nor02ii port map ( Y=>nx2790, A0=>nx28856, A1=>nx36105);
   ix2785 : xor2 port map ( Y=>nx12975, A0=>nx28873, A1=>nx29024);
   ix2773 : xor2 port map ( Y=>nx12977, A0=>nx28903, A1=>nx35417);
   ix15264 : mux21_ni port map ( Y=>nx15263, A0=>
      booth_booth_integrtaion_2_booth_output_24, A1=>nx2766, S0=>nx36099);
   ix2767 : nor02ii port map ( Y=>nx2766, A0=>nx28891, A1=>nx36107);
   ix2761 : xor2 port map ( Y=>nx12978, A0=>nx28908, A1=>nx29021);
   ix2749 : xor2 port map ( Y=>nx12979, A0=>nx28938, A1=>nx35419);
   ix15244 : mux21_ni port map ( Y=>nx15243, A0=>
      booth_booth_integrtaion_2_booth_output_26, A1=>nx2742, S0=>nx36099);
   ix2743 : nor02ii port map ( Y=>nx2742, A0=>nx28926, A1=>nx36107);
   ix2737 : xor2 port map ( Y=>nx12981, A0=>nx28943, A1=>nx29018);
   ix2725 : xor2 port map ( Y=>nx12983, A0=>nx28973, A1=>nx35421);
   ix15224 : mux21_ni port map ( Y=>nx15223, A0=>
      booth_booth_integrtaion_2_booth_output_28, A1=>nx2718, S0=>nx35403);
   ix2719 : nor02ii port map ( Y=>nx2718, A0=>nx28961, A1=>nx36107);
   ix2713 : xor2 port map ( Y=>nx12985, A0=>nx28978, A1=>nx29015);
   ix2701 : xor2 port map ( Y=>nx12987, A0=>nx29008, A1=>nx35423);
   ix15204 : mux21_ni port map ( Y=>nx15203, A0=>
      booth_booth_integrtaion_2_booth_output_31, A1=>nx2694, S0=>nx35403);
   ix2695 : nor02ii port map ( Y=>nx2694, A0=>nx28996, A1=>nx36107);
   ix2689 : xor2 port map ( Y=>nx2688, A0=>nx29008, A1=>nx29011);
   ix2875 : nor02ii port map ( Y=>nx2874, A0=>nx2338, A1=>nx36107);
   ix24264 : ao32 port map ( Y=>nx24263, A0=>nx35959, A1=>nx35645, A2=>
      nx36291, B0=>max_calc_ans3_0, B1=>nx35877);
   ix29058 : mux21 port map ( Y=>nx35645, A0=>nx29502, A1=>nx29061, S0=>
      nx35887);
   ix20194 : mux21_ni port map ( Y=>nx20193, A0=>label_5_output(0), A1=>
      label_5_input_0, S0=>nx36251);
   ix20184 : mux21_ni port map ( Y=>nx20183, A0=>
      label_5_input_state_machine_0, A1=>mdr_data_out(64), S0=>nx36211);
   ix20174 : mux21_ni port map ( Y=>nx20173, A0=>nx35763, A1=>nx10374, S0=>
      nx35431);
   ix10375 : mux21_ni port map ( Y=>nx10374, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_4_1, S0=>nx36117);
   ix20164 : mux21_ni port map ( Y=>nx20163, A0=>
      booth_booth_integration_output_4_1, A1=>nx10362, S0=>nx35431);
   ix10363 : mux21_ni port map ( Y=>nx10362, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_4_2, S0=>nx36117);
   ix20154 : mux21_ni port map ( Y=>nx20153, A0=>
      booth_booth_integration_output_4_2, A1=>nx10350, S0=>nx35431);
   ix10351 : mux21_ni port map ( Y=>nx10350, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_4_3, S0=>nx36117);
   ix20144 : mux21_ni port map ( Y=>nx20143, A0=>
      booth_booth_integration_output_4_3, A1=>nx10338, S0=>nx35431);
   ix10339 : mux21_ni port map ( Y=>nx10338, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_4_4, S0=>nx36117);
   ix20134 : mux21_ni port map ( Y=>nx20133, A0=>
      booth_booth_integration_output_4_4, A1=>nx10326, S0=>nx35431);
   ix10327 : mux21_ni port map ( Y=>nx10326, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_4_5, S0=>nx36117);
   ix20124 : mux21_ni port map ( Y=>nx20123, A0=>
      booth_booth_integration_output_4_5, A1=>nx10314, S0=>nx35431);
   ix10315 : mux21_ni port map ( Y=>nx10314, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_4_6, S0=>nx36119);
   ix20114 : mux21_ni port map ( Y=>nx20113, A0=>
      booth_booth_integration_output_4_6, A1=>nx10302, S0=>nx35431);
   ix10303 : mux21_ni port map ( Y=>nx10302, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_4_7, S0=>nx36119);
   ix20104 : mux21_ni port map ( Y=>nx20103, A0=>
      booth_booth_integration_output_4_7, A1=>nx10290, S0=>nx36109);
   ix10291 : mux21_ni port map ( Y=>nx10290, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_4_8, S0=>nx36119);
   ix20094 : mux21_ni port map ( Y=>nx20093, A0=>
      booth_booth_integration_output_4_8, A1=>nx10278, S0=>nx36109);
   ix10279 : mux21_ni port map ( Y=>nx10278, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_4_9, S0=>nx36119);
   ix20084 : mux21_ni port map ( Y=>nx20083, A0=>
      booth_booth_integration_output_4_9, A1=>nx10266, S0=>nx36109);
   ix10267 : mux21_ni port map ( Y=>nx10266, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_4_10, S0=>nx36119);
   ix20074 : mux21_ni port map ( Y=>nx20073, A0=>
      booth_booth_integration_output_4_10, A1=>nx10254, S0=>nx36111);
   ix10255 : mux21_ni port map ( Y=>nx10254, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_4_11, S0=>nx36119);
   ix20064 : mux21_ni port map ( Y=>nx20063, A0=>
      booth_booth_integration_output_4_11, A1=>nx10242, S0=>nx36111);
   ix10243 : mux21_ni port map ( Y=>nx10242, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_4_12, S0=>nx36119);
   ix20054 : mux21_ni port map ( Y=>nx20053, A0=>
      booth_booth_integration_output_4_12, A1=>nx10230, S0=>nx36111);
   ix10231 : mux21_ni port map ( Y=>nx10230, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_4_13, S0=>nx36121);
   ix20044 : mux21_ni port map ( Y=>nx20043, A0=>
      booth_booth_integration_output_4_13, A1=>nx10218, S0=>nx36111);
   ix10219 : mux21_ni port map ( Y=>nx10218, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_4_14, S0=>nx36121);
   ix20034 : mux21_ni port map ( Y=>nx20033, A0=>
      booth_booth_integration_output_4_14, A1=>nx10206, S0=>nx36111);
   ix10207 : mux21_ni port map ( Y=>nx10206, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_4_15, S0=>nx36121);
   ix20024 : mux21 port map ( Y=>nx20023, A0=>nx29480, A1=>nx29122, S0=>
      nx36111);
   ix19674 : mux21_ni port map ( Y=>nx19673, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_0, A1=>nx34939, S0=>nx35823
   );
   ix19660 : and02 port map ( Y=>nx19659, A0=>nx36349, A1=>
      booth_booth_integrtaion_4_shift_Reg_count_0);
   ix19854 : mux21_ni port map ( Y=>nx19853, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_9, A1=>nx34925, S0=>nx35823
   );
   ix19844 : mux21_ni port map ( Y=>nx19843, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_8, S0=>nx36111);
   ix19834 : mux21_ni port map ( Y=>nx19833, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_8, S0=>nx35823);
   ix19824 : mux21_ni port map ( Y=>nx19823, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_7, S0=>nx36113);
   ix19814 : mux21_ni port map ( Y=>nx19813, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_7, S0=>nx35823);
   ix19804 : mux21_ni port map ( Y=>nx19803, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_6, S0=>nx36113);
   ix19794 : mux21_ni port map ( Y=>nx19793, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_6, S0=>nx35823);
   ix19784 : mux21_ni port map ( Y=>nx19783, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_5, S0=>nx36113);
   ix19774 : mux21_ni port map ( Y=>nx19773, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_5, S0=>nx35823);
   ix19764 : mux21_ni port map ( Y=>nx19763, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_4, S0=>nx36113);
   ix19754 : mux21_ni port map ( Y=>nx19753, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_4, S0=>nx35825);
   ix19744 : mux21_ni port map ( Y=>nx19743, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_3, S0=>nx36113);
   ix19734 : mux21_ni port map ( Y=>nx19733, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_3, S0=>nx35825);
   ix19724 : mux21_ni port map ( Y=>nx19723, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_2, S0=>nx36113);
   ix19714 : mux21_ni port map ( Y=>nx19713, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_2, S0=>nx35825);
   ix19704 : mux21_ni port map ( Y=>nx19703, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_1, S0=>nx36113);
   ix19694 : mux21_ni port map ( Y=>nx19693, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_4_shift_Reg_output_1, S0=>nx35825);
   ix19684 : mux21_ni port map ( Y=>nx19683, A0=>
      booth_booth_integrtaion_4_shift_Reg_count_1, A1=>nx34939, S0=>nx36115
   );
   ix9647 : and02 port map ( Y=>nx9646, A0=>nx29195, A1=>nx35763);
   ix29198 : or03 port map ( Y=>nx29197, A0=>nx29199, A1=>
      booth_booth_integrtaion_4_shift_reg_output_0, A2=>nx36349);
   ix20014 : mux21_ni port map ( Y=>nx20013, A0=>
      booth_booth_integrtaion_4_booth_output_16, A1=>nx10176, S0=>nx36115);
   ix10177 : nor02ii port map ( Y=>nx10176, A0=>nx29206, A1=>nx36121);
   ix9653 : nor02ii port map ( Y=>nx9652, A0=>nx29190, A1=>
      booth_booth_integrtaion_4_booth_output_16);
   ix10171 : xor2 port map ( Y=>nx13217, A0=>nx29212, A1=>nx29476);
   ix10159 : xor2 port map ( Y=>nx13219, A0=>nx29237, A1=>nx35437);
   ix19994 : mux21_ni port map ( Y=>nx19993, A0=>
      booth_booth_integrtaion_4_booth_output_18, A1=>nx10152, S0=>nx36115);
   ix10153 : nor02ii port map ( Y=>nx10152, A0=>nx29227, A1=>nx36121);
   ix10147 : xor2 port map ( Y=>nx13221, A0=>nx29242, A1=>nx29473);
   ix29259 : or02 port map ( Y=>nx29258, A0=>nx29195, A1=>nx35765);
   ix10135 : xor2 port map ( Y=>nx13223, A0=>nx29276, A1=>nx35439);
   ix19974 : mux21_ni port map ( Y=>nx19973, A0=>
      booth_booth_integrtaion_4_booth_output_20, A1=>nx10128, S0=>nx36115);
   ix10129 : nor02ii port map ( Y=>nx10128, A0=>nx29264, A1=>nx36121);
   ix10123 : xor2 port map ( Y=>nx13224, A0=>nx29281, A1=>nx29470);
   ix10111 : xor2 port map ( Y=>nx13225, A0=>nx29311, A1=>nx35441);
   ix19954 : mux21_ni port map ( Y=>nx19953, A0=>
      booth_booth_integrtaion_4_booth_output_22, A1=>nx10104, S0=>nx36115);
   ix10105 : nor02ii port map ( Y=>nx10104, A0=>nx29299, A1=>nx36121);
   ix10099 : xor2 port map ( Y=>nx13226, A0=>nx29316, A1=>nx29467);
   ix10087 : xor2 port map ( Y=>nx13227, A0=>nx29346, A1=>nx35443);
   ix19934 : mux21_ni port map ( Y=>nx19933, A0=>
      booth_booth_integrtaion_4_booth_output_24, A1=>nx10080, S0=>nx36115);
   ix10081 : nor02ii port map ( Y=>nx10080, A0=>nx29334, A1=>nx36123);
   ix10075 : xor2 port map ( Y=>nx13228, A0=>nx29351, A1=>nx29464);
   ix10063 : xor2 port map ( Y=>nx13229, A0=>nx29381, A1=>nx35445);
   ix19914 : mux21_ni port map ( Y=>nx19913, A0=>
      booth_booth_integrtaion_4_booth_output_26, A1=>nx10056, S0=>nx36115);
   ix10057 : nor02ii port map ( Y=>nx10056, A0=>nx29369, A1=>nx36123);
   ix10051 : xor2 port map ( Y=>nx13231, A0=>nx29386, A1=>nx29461);
   ix10039 : xor2 port map ( Y=>nx13233, A0=>nx29416, A1=>nx35447);
   ix19894 : mux21_ni port map ( Y=>nx19893, A0=>
      booth_booth_integrtaion_4_booth_output_28, A1=>nx10032, S0=>nx35429);
   ix10033 : nor02ii port map ( Y=>nx10032, A0=>nx29404, A1=>nx36123);
   ix10027 : xor2 port map ( Y=>nx13235, A0=>nx29421, A1=>nx29458);
   ix10015 : xor2 port map ( Y=>nx13236, A0=>nx29451, A1=>nx35449);
   ix19874 : mux21_ni port map ( Y=>nx19873, A0=>
      booth_booth_integrtaion_4_booth_output_31, A1=>nx10008, S0=>nx35429);
   ix10009 : nor02ii port map ( Y=>nx10008, A0=>nx29439, A1=>nx36123);
   ix10003 : xor2 port map ( Y=>nx10002, A0=>nx29451, A1=>nx29454);
   ix10189 : nor02ii port map ( Y=>nx10188, A0=>nx9652, A1=>nx36123);
   ix29499 : and04 port map ( Y=>nx29498, A0=>max_calc_state_0, A1=>nx35979, 
      A2=>nx35959, A3=>nx26203);
   ix21034 : mux21_ni port map ( Y=>nx21033, A0=>label_6_output(0), A1=>
      label_6_input_0, S0=>nx36251);
   ix21024 : mux21_ni port map ( Y=>nx21023, A0=>
      label_6_input_state_machine_0, A1=>mdr_data_out(80), S0=>nx36211);
   ix21014 : mux21_ni port map ( Y=>nx21013, A0=>nx35767, A1=>nx11696, S0=>
      nx35479);
   ix11697 : mux21_ni port map ( Y=>nx11696, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_5_1, S0=>nx36139);
   ix21004 : mux21_ni port map ( Y=>nx21003, A0=>
      booth_booth_integration_output_5_1, A1=>nx11684, S0=>nx35479);
   ix11685 : mux21_ni port map ( Y=>nx11684, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_5_2, S0=>nx36139);
   ix20994 : mux21_ni port map ( Y=>nx20993, A0=>
      booth_booth_integration_output_5_2, A1=>nx11672, S0=>nx35479);
   ix11673 : mux21_ni port map ( Y=>nx11672, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_5_3, S0=>nx36139);
   ix20984 : mux21_ni port map ( Y=>nx20983, A0=>
      booth_booth_integration_output_5_3, A1=>nx11660, S0=>nx35479);
   ix11661 : mux21_ni port map ( Y=>nx11660, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_5_4, S0=>nx36139);
   ix20974 : mux21_ni port map ( Y=>nx20973, A0=>
      booth_booth_integration_output_5_4, A1=>nx11648, S0=>nx35479);
   ix11649 : mux21_ni port map ( Y=>nx11648, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_5_5, S0=>nx36139);
   ix20964 : mux21_ni port map ( Y=>nx20963, A0=>
      booth_booth_integration_output_5_5, A1=>nx11636, S0=>nx35479);
   ix11637 : mux21_ni port map ( Y=>nx11636, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_5_6, S0=>nx36141);
   ix20954 : mux21_ni port map ( Y=>nx20953, A0=>
      booth_booth_integration_output_5_6, A1=>nx11624, S0=>nx35479);
   ix11625 : mux21_ni port map ( Y=>nx11624, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_5_7, S0=>nx36141);
   ix20944 : mux21_ni port map ( Y=>nx20943, A0=>
      booth_booth_integration_output_5_7, A1=>nx11612, S0=>nx36131);
   ix11613 : mux21_ni port map ( Y=>nx11612, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_5_8, S0=>nx36141);
   ix20934 : mux21_ni port map ( Y=>nx20933, A0=>
      booth_booth_integration_output_5_8, A1=>nx11600, S0=>nx36131);
   ix11601 : mux21_ni port map ( Y=>nx11600, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_5_9, S0=>nx36141);
   ix20924 : mux21_ni port map ( Y=>nx20923, A0=>
      booth_booth_integration_output_5_9, A1=>nx11588, S0=>nx36131);
   ix11589 : mux21_ni port map ( Y=>nx11588, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_5_10, S0=>nx36141);
   ix20914 : mux21_ni port map ( Y=>nx20913, A0=>
      booth_booth_integration_output_5_10, A1=>nx11576, S0=>nx36133);
   ix11577 : mux21_ni port map ( Y=>nx11576, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_5_11, S0=>nx36141);
   ix20904 : mux21_ni port map ( Y=>nx20903, A0=>
      booth_booth_integration_output_5_11, A1=>nx11564, S0=>nx36133);
   ix11565 : mux21_ni port map ( Y=>nx11564, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_5_12, S0=>nx36141);
   ix20894 : mux21_ni port map ( Y=>nx20893, A0=>
      booth_booth_integration_output_5_12, A1=>nx11552, S0=>nx36133);
   ix11553 : mux21_ni port map ( Y=>nx11552, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_5_13, S0=>nx36143);
   ix20884 : mux21_ni port map ( Y=>nx20883, A0=>
      booth_booth_integration_output_5_13, A1=>nx11540, S0=>nx36133);
   ix11541 : mux21_ni port map ( Y=>nx11540, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_5_14, S0=>nx36143);
   ix20874 : mux21_ni port map ( Y=>nx20873, A0=>
      booth_booth_integration_output_5_14, A1=>nx11528, S0=>nx36133);
   ix11529 : mux21_ni port map ( Y=>nx11528, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_5_15, S0=>nx36143);
   ix20864 : mux21 port map ( Y=>nx20863, A0=>nx29921, A1=>nx29563, S0=>
      nx36133);
   ix20514 : mux21_ni port map ( Y=>nx20513, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_0, A1=>nx34971, S0=>nx35827
   );
   ix20500 : and02 port map ( Y=>nx20499, A0=>nx36353, A1=>
      booth_booth_integrtaion_5_shift_Reg_count_0);
   ix20694 : mux21_ni port map ( Y=>nx20693, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_9, A1=>nx34957, S0=>nx35827
   );
   ix20684 : mux21_ni port map ( Y=>nx20683, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_8, S0=>nx36133);
   ix20674 : mux21_ni port map ( Y=>nx20673, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_8, S0=>nx35827);
   ix20664 : mux21_ni port map ( Y=>nx20663, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_7, S0=>nx36135);
   ix20654 : mux21_ni port map ( Y=>nx20653, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_7, S0=>nx35827);
   ix20644 : mux21_ni port map ( Y=>nx20643, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_6, S0=>nx36135);
   ix20634 : mux21_ni port map ( Y=>nx20633, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_6, S0=>nx35827);
   ix20624 : mux21_ni port map ( Y=>nx20623, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_5, S0=>nx36135);
   ix20614 : mux21_ni port map ( Y=>nx20613, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_5, S0=>nx35827);
   ix20604 : mux21_ni port map ( Y=>nx20603, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_4, S0=>nx36135);
   ix20594 : mux21_ni port map ( Y=>nx20593, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_4, S0=>nx35829);
   ix20584 : mux21_ni port map ( Y=>nx20583, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_3, S0=>nx36135);
   ix20574 : mux21_ni port map ( Y=>nx20573, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_3, S0=>nx35829);
   ix20564 : mux21_ni port map ( Y=>nx20563, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_2, S0=>nx36135);
   ix20554 : mux21_ni port map ( Y=>nx20553, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_2, S0=>nx35829);
   ix20544 : mux21_ni port map ( Y=>nx20543, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_1, S0=>nx36135);
   ix20534 : mux21_ni port map ( Y=>nx20533, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_5_shift_Reg_output_1, S0=>nx35829);
   ix20524 : mux21_ni port map ( Y=>nx20523, A0=>
      booth_booth_integrtaion_5_shift_Reg_count_1, A1=>nx34971, S0=>nx36137
   );
   ix10969 : and02 port map ( Y=>nx10968, A0=>nx29636, A1=>nx35767);
   ix29639 : or03 port map ( Y=>nx29638, A0=>nx29640, A1=>
      booth_booth_integrtaion_5_shift_reg_output_0, A2=>nx36353);
   ix20854 : mux21_ni port map ( Y=>nx20853, A0=>
      booth_booth_integrtaion_5_booth_output_16, A1=>nx11498, S0=>nx36137);
   ix11499 : nor02ii port map ( Y=>nx11498, A0=>nx29647, A1=>nx36143);
   ix10975 : nor02ii port map ( Y=>nx10974, A0=>nx29631, A1=>
      booth_booth_integrtaion_5_booth_output_16);
   ix11493 : xor2 port map ( Y=>nx13257, A0=>nx29653, A1=>nx29917);
   ix11481 : xor2 port map ( Y=>nx13259, A0=>nx29678, A1=>nx35485);
   ix20834 : mux21_ni port map ( Y=>nx20833, A0=>
      booth_booth_integrtaion_5_booth_output_18, A1=>nx11474, S0=>nx36137);
   ix11475 : nor02ii port map ( Y=>nx11474, A0=>nx29668, A1=>nx36143);
   ix11469 : xor2 port map ( Y=>nx13260, A0=>nx29683, A1=>nx29914);
   ix29700 : or02 port map ( Y=>nx29699, A0=>nx29636, A1=>nx35769);
   ix11457 : xor2 port map ( Y=>nx13261, A0=>nx29717, A1=>nx35487);
   ix20814 : mux21_ni port map ( Y=>nx20813, A0=>
      booth_booth_integrtaion_5_booth_output_20, A1=>nx11450, S0=>nx36137);
   ix11451 : nor02ii port map ( Y=>nx11450, A0=>nx29705, A1=>nx36143);
   ix11445 : xor2 port map ( Y=>nx13262, A0=>nx29722, A1=>nx29911);
   ix11433 : xor2 port map ( Y=>nx13263, A0=>nx29752, A1=>nx35489);
   ix20794 : mux21_ni port map ( Y=>nx20793, A0=>
      booth_booth_integrtaion_5_booth_output_22, A1=>nx11426, S0=>nx36137);
   ix11427 : nor02ii port map ( Y=>nx11426, A0=>nx29740, A1=>nx36143);
   ix11421 : xor2 port map ( Y=>nx13264, A0=>nx29757, A1=>nx29908);
   ix11409 : xor2 port map ( Y=>nx13265, A0=>nx29787, A1=>nx35491);
   ix20774 : mux21_ni port map ( Y=>nx20773, A0=>
      booth_booth_integrtaion_5_booth_output_24, A1=>nx11402, S0=>nx36137);
   ix11403 : nor02ii port map ( Y=>nx11402, A0=>nx29775, A1=>nx36145);
   ix11397 : xor2 port map ( Y=>nx13267, A0=>nx29792, A1=>nx29905);
   ix11385 : xor2 port map ( Y=>nx13269, A0=>nx29822, A1=>nx35493);
   ix20754 : mux21_ni port map ( Y=>nx20753, A0=>
      booth_booth_integrtaion_5_booth_output_26, A1=>nx11378, S0=>nx36137);
   ix11379 : nor02ii port map ( Y=>nx11378, A0=>nx29810, A1=>nx36145);
   ix11373 : xor2 port map ( Y=>nx13271, A0=>nx29827, A1=>nx29902);
   ix11361 : xor2 port map ( Y=>nx13272, A0=>nx29857, A1=>nx35495);
   ix20734 : mux21_ni port map ( Y=>nx20733, A0=>
      booth_booth_integrtaion_5_booth_output_28, A1=>nx11354, S0=>nx35477);
   ix11355 : nor02ii port map ( Y=>nx11354, A0=>nx29845, A1=>nx36145);
   ix11349 : xor2 port map ( Y=>nx13273, A0=>nx29862, A1=>nx29899);
   ix11337 : xor2 port map ( Y=>nx13274, A0=>nx29892, A1=>nx35497);
   ix20714 : mux21_ni port map ( Y=>nx20713, A0=>
      booth_booth_integrtaion_5_booth_output_31, A1=>nx11330, S0=>nx35477);
   ix11331 : nor02ii port map ( Y=>nx11330, A0=>nx29880, A1=>nx36145);
   ix11325 : xor2 port map ( Y=>nx11324, A0=>nx29892, A1=>nx29895);
   ix11511 : nor02ii port map ( Y=>nx11510, A0=>nx10974, A1=>nx36145);
   ix29946 : or03 port map ( Y=>nx29945, A0=>nx30129, A1=>nx36195, A2=>
      nx36069);
   ix21304 : mux21_ni port map ( Y=>nx21303, A0=>label_6_output(14), A1=>
      label_6_input_14, S0=>nx36253);
   ix12155 : mux21_ni port map ( Y=>nx12154, A0=>nx12150, A1=>
      label_6_input_state_machine_14, S0=>nx35927);
   ix20484 : mux21_ni port map ( Y=>nx20483, A0=>
      label_6_input_state_machine_14, A1=>mdr_data_out(94), S0=>nx36211);
   ix21294 : mux21_ni port map ( Y=>nx21293, A0=>label_6_output(13), A1=>
      label_6_input_13, S0=>nx36253);
   ix12129 : mux21_ni port map ( Y=>nx12128, A0=>nx12124, A1=>
      label_6_input_state_machine_13, S0=>nx35927);
   ix21284 : mux21_ni port map ( Y=>nx21283, A0=>
      label_6_input_state_machine_13, A1=>mdr_data_out(93), S0=>nx36211);
   ix21254 : mux21_ni port map ( Y=>nx21253, A0=>label_6_output(11), A1=>
      label_6_input_11, S0=>nx36251);
   ix12065 : mux21_ni port map ( Y=>nx12064, A0=>nx12060, A1=>
      label_6_input_state_machine_11, S0=>nx35927);
   ix21244 : mux21_ni port map ( Y=>nx21243, A0=>
      label_6_input_state_machine_11, A1=>mdr_data_out(91), S0=>nx36211);
   ix21214 : mux21_ni port map ( Y=>nx21213, A0=>label_6_output(9), A1=>
      label_6_input_9, S0=>nx36251);
   ix12001 : mux21_ni port map ( Y=>nx12000, A0=>nx11996, A1=>
      label_6_input_state_machine_9, S0=>nx35927);
   ix21204 : mux21_ni port map ( Y=>nx21203, A0=>
      label_6_input_state_machine_9, A1=>mdr_data_out(89), S0=>nx35595);
   ix21174 : mux21_ni port map ( Y=>nx21173, A0=>label_6_output(7), A1=>
      label_6_input_7, S0=>nx36251);
   ix11937 : mux21_ni port map ( Y=>nx11936, A0=>nx11932, A1=>
      label_6_input_state_machine_7, S0=>nx35929);
   ix21164 : mux21_ni port map ( Y=>nx21163, A0=>
      label_6_input_state_machine_7, A1=>mdr_data_out(87), S0=>nx36213);
   ix21134 : mux21_ni port map ( Y=>nx21133, A0=>label_6_output(5), A1=>
      label_6_input_5, S0=>nx36251);
   ix11873 : mux21_ni port map ( Y=>nx11872, A0=>nx11868, A1=>
      label_6_input_state_machine_5, S0=>nx35929);
   ix21124 : mux21_ni port map ( Y=>nx21123, A0=>
      label_6_input_state_machine_5, A1=>mdr_data_out(85), S0=>nx36213);
   ix21094 : mux21_ni port map ( Y=>nx21093, A0=>label_6_output(3), A1=>
      label_6_input_3, S0=>nx36251);
   ix11809 : mux21_ni port map ( Y=>nx11808, A0=>nx11804, A1=>
      label_6_input_state_machine_3, S0=>nx35929);
   ix21084 : mux21_ni port map ( Y=>nx21083, A0=>
      label_6_input_state_machine_3, A1=>mdr_data_out(83), S0=>nx36213);
   ix21054 : mux21_ni port map ( Y=>nx21053, A0=>label_6_output(1), A1=>
      label_6_input_1, S0=>nx36391);
   ix11745 : mux21_ni port map ( Y=>nx11744, A0=>nx11740, A1=>
      label_6_input_state_machine_1, S0=>nx35929);
   ix21044 : mux21_ni port map ( Y=>nx21043, A0=>
      label_6_input_state_machine_1, A1=>mdr_data_out(81), S0=>nx36213);
   ix30038 : xnor2 port map ( Y=>nx30037, A0=>nx29935, A1=>nx30047);
   ix21074 : mux21_ni port map ( Y=>nx21073, A0=>label_6_output(2), A1=>
      label_6_input_2, S0=>nx36391);
   ix11777 : mux21_ni port map ( Y=>nx11776, A0=>nx11772, A1=>
      label_6_input_state_machine_2, S0=>nx35929);
   ix21064 : mux21_ni port map ( Y=>nx21063, A0=>
      label_6_input_state_machine_2, A1=>mdr_data_out(82), S0=>nx36213);
   ix30053 : xnor2 port map ( Y=>nx30052, A0=>nx29933, A1=>nx30062);
   ix21114 : mux21_ni port map ( Y=>nx21113, A0=>label_6_output(4), A1=>
      label_6_input_4, S0=>nx36391);
   ix11841 : mux21_ni port map ( Y=>nx11840, A0=>nx11836, A1=>
      label_6_input_state_machine_4, S0=>nx35929);
   ix21104 : mux21_ni port map ( Y=>nx21103, A0=>
      label_6_input_state_machine_4, A1=>mdr_data_out(84), S0=>nx36213);
   ix30068 : xnor2 port map ( Y=>nx30067, A0=>nx29931, A1=>nx30077);
   ix21154 : mux21_ni port map ( Y=>nx21153, A0=>label_6_output(6), A1=>
      label_6_input_6, S0=>nx36391);
   ix11905 : mux21_ni port map ( Y=>nx11904, A0=>nx11900, A1=>
      label_6_input_state_machine_6, S0=>nx35929);
   ix21144 : mux21_ni port map ( Y=>nx21143, A0=>
      label_6_input_state_machine_6, A1=>mdr_data_out(86), S0=>nx36213);
   ix30083 : xnor2 port map ( Y=>nx30082, A0=>nx29929, A1=>nx30092);
   ix21194 : mux21_ni port map ( Y=>nx21193, A0=>label_6_output(8), A1=>
      label_6_input_8, S0=>nx36391);
   ix11969 : mux21_ni port map ( Y=>nx11968, A0=>nx11964, A1=>
      label_6_input_state_machine_8, S0=>nx35931);
   ix21184 : mux21_ni port map ( Y=>nx21183, A0=>
      label_6_input_state_machine_8, A1=>mdr_data_out(88), S0=>nx36215);
   ix30098 : xnor2 port map ( Y=>nx30097, A0=>nx29927, A1=>nx30107);
   ix21234 : mux21_ni port map ( Y=>nx21233, A0=>label_6_output(10), A1=>
      label_6_input_10, S0=>nx36391);
   ix12033 : mux21_ni port map ( Y=>nx12032, A0=>nx12028, A1=>
      label_6_input_state_machine_10, S0=>nx35931);
   ix21224 : mux21_ni port map ( Y=>nx21223, A0=>
      label_6_input_state_machine_10, A1=>mdr_data_out(90), S0=>nx36215);
   ix30113 : xnor2 port map ( Y=>nx30112, A0=>nx29925, A1=>nx30122);
   ix21274 : mux21_ni port map ( Y=>nx21273, A0=>label_6_output(12), A1=>
      label_6_input_12, S0=>nx36391);
   ix12097 : mux21_ni port map ( Y=>nx12096, A0=>nx12092, A1=>
      label_6_input_state_machine_12, S0=>nx35931);
   ix21264 : mux21_ni port map ( Y=>nx21263, A0=>
      label_6_input_state_machine_12, A1=>mdr_data_out(92), S0=>nx36215);
   ix30128 : xnor2 port map ( Y=>nx30127, A0=>nx29923, A1=>nx30129);
   ix30135 : or03 port map ( Y=>nx30134, A0=>nx30318, A1=>nx36195, A2=>
      nx36069);
   ix20464 : mux21_ni port map ( Y=>nx20463, A0=>label_5_output(14), A1=>
      label_5_input_14, S0=>nx36253);
   ix10833 : mux21_ni port map ( Y=>nx10832, A0=>nx10828, A1=>
      label_5_input_state_machine_14, S0=>nx35931);
   ix19644 : mux21_ni port map ( Y=>nx19643, A0=>
      label_5_input_state_machine_14, A1=>mdr_data_out(78), S0=>nx36215);
   ix20454 : mux21_ni port map ( Y=>nx20453, A0=>label_5_output(13), A1=>
      label_5_input_13, S0=>nx36253);
   ix10807 : mux21_ni port map ( Y=>nx10806, A0=>nx10802, A1=>
      label_5_input_state_machine_13, S0=>nx35931);
   ix20444 : mux21_ni port map ( Y=>nx20443, A0=>
      label_5_input_state_machine_13, A1=>mdr_data_out(77), S0=>nx36215);
   ix20414 : mux21_ni port map ( Y=>nx20413, A0=>label_5_output(11), A1=>
      label_5_input_11, S0=>nx36253);
   ix10743 : mux21_ni port map ( Y=>nx10742, A0=>nx10738, A1=>
      label_5_input_state_machine_11, S0=>nx35931);
   ix20404 : mux21_ni port map ( Y=>nx20403, A0=>
      label_5_input_state_machine_11, A1=>mdr_data_out(75), S0=>nx36215);
   ix20374 : mux21_ni port map ( Y=>nx20373, A0=>label_5_output(9), A1=>
      label_5_input_9, S0=>nx36253);
   ix10679 : mux21_ni port map ( Y=>nx10678, A0=>nx10674, A1=>
      label_5_input_state_machine_9, S0=>nx35931);
   ix20364 : mux21_ni port map ( Y=>nx20363, A0=>
      label_5_input_state_machine_9, A1=>mdr_data_out(73), S0=>nx36215);
   ix20334 : mux21_ni port map ( Y=>nx20333, A0=>label_5_output(7), A1=>
      label_5_input_7, S0=>nx36253);
   ix10615 : mux21_ni port map ( Y=>nx10614, A0=>nx10610, A1=>
      label_5_input_state_machine_7, S0=>nx35933);
   ix20324 : mux21_ni port map ( Y=>nx20323, A0=>
      label_5_input_state_machine_7, A1=>mdr_data_out(71), S0=>nx36217);
   ix20294 : mux21_ni port map ( Y=>nx20293, A0=>label_5_output(5), A1=>
      label_5_input_5, S0=>nx36255);
   ix10551 : mux21_ni port map ( Y=>nx10550, A0=>nx10546, A1=>
      label_5_input_state_machine_5, S0=>nx35933);
   ix20284 : mux21_ni port map ( Y=>nx20283, A0=>
      label_5_input_state_machine_5, A1=>mdr_data_out(69), S0=>nx36217);
   ix20254 : mux21_ni port map ( Y=>nx20253, A0=>label_5_output(3), A1=>
      label_5_input_3, S0=>nx36255);
   ix10487 : mux21_ni port map ( Y=>nx10486, A0=>nx10482, A1=>
      label_5_input_state_machine_3, S0=>nx35933);
   ix20244 : mux21_ni port map ( Y=>nx20243, A0=>
      label_5_input_state_machine_3, A1=>mdr_data_out(67), S0=>nx36217);
   ix20214 : mux21_ni port map ( Y=>nx20213, A0=>label_5_output(1), A1=>
      label_5_input_1, S0=>nx36255);
   ix10423 : mux21_ni port map ( Y=>nx10422, A0=>nx10418, A1=>
      label_5_input_state_machine_1, S0=>nx35933);
   ix20204 : mux21_ni port map ( Y=>nx20203, A0=>
      label_5_input_state_machine_1, A1=>mdr_data_out(65), S0=>nx36217);
   ix30227 : xnor2 port map ( Y=>nx30226, A0=>nx29494, A1=>nx30236);
   ix20234 : mux21_ni port map ( Y=>nx20233, A0=>label_5_output(2), A1=>
      label_5_input_2, S0=>nx36255);
   ix10455 : mux21_ni port map ( Y=>nx10454, A0=>nx10450, A1=>
      label_5_input_state_machine_2, S0=>nx35933);
   ix20224 : mux21_ni port map ( Y=>nx20223, A0=>
      label_5_input_state_machine_2, A1=>mdr_data_out(66), S0=>nx36217);
   ix30242 : xnor2 port map ( Y=>nx30241, A0=>nx29492, A1=>nx30251);
   ix20274 : mux21_ni port map ( Y=>nx20273, A0=>label_5_output(4), A1=>
      label_5_input_4, S0=>nx36255);
   ix10519 : mux21_ni port map ( Y=>nx10518, A0=>nx10514, A1=>
      label_5_input_state_machine_4, S0=>nx35933);
   ix20264 : mux21_ni port map ( Y=>nx20263, A0=>
      label_5_input_state_machine_4, A1=>mdr_data_out(68), S0=>nx36217);
   ix30257 : xnor2 port map ( Y=>nx30256, A0=>nx29490, A1=>nx30266);
   ix20314 : mux21_ni port map ( Y=>nx20313, A0=>label_5_output(6), A1=>
      label_5_input_6, S0=>nx36255);
   ix10583 : mux21_ni port map ( Y=>nx10582, A0=>nx10578, A1=>
      label_5_input_state_machine_6, S0=>nx35933);
   ix20304 : mux21_ni port map ( Y=>nx20303, A0=>
      label_5_input_state_machine_6, A1=>mdr_data_out(70), S0=>nx36217);
   ix30272 : xnor2 port map ( Y=>nx30271, A0=>nx29488, A1=>nx30281);
   ix20354 : mux21_ni port map ( Y=>nx20353, A0=>label_5_output(8), A1=>
      label_5_input_8, S0=>nx36255);
   ix10647 : mux21_ni port map ( Y=>nx10646, A0=>nx10642, A1=>
      label_5_input_state_machine_8, S0=>nx35935);
   ix20344 : mux21_ni port map ( Y=>nx20343, A0=>
      label_5_input_state_machine_8, A1=>mdr_data_out(72), S0=>nx36219);
   ix30287 : xnor2 port map ( Y=>nx30286, A0=>nx29486, A1=>nx30296);
   ix20394 : mux21_ni port map ( Y=>nx20393, A0=>label_5_output(10), A1=>
      label_5_input_10, S0=>nx36257);
   ix10711 : mux21_ni port map ( Y=>nx10710, A0=>nx10706, A1=>
      label_5_input_state_machine_10, S0=>nx35935);
   ix20384 : mux21_ni port map ( Y=>nx20383, A0=>
      label_5_input_state_machine_10, A1=>mdr_data_out(74), S0=>nx36219);
   ix30302 : xnor2 port map ( Y=>nx30301, A0=>nx29484, A1=>nx30311);
   ix20434 : mux21_ni port map ( Y=>nx20433, A0=>label_5_output(12), A1=>
      label_5_input_12, S0=>nx36257);
   ix10775 : mux21_ni port map ( Y=>nx10774, A0=>nx10770, A1=>
      label_5_input_state_machine_12, S0=>nx35935);
   ix20424 : mux21_ni port map ( Y=>nx20423, A0=>
      label_5_input_state_machine_12, A1=>mdr_data_out(76), S0=>nx36219);
   ix30317 : xnor2 port map ( Y=>nx30316, A0=>nx29482, A1=>nx30318);
   ix12177 : xnor2 port map ( Y=>nx12176, A0=>nx29942, A1=>nx30132);
   ix30322 : xnor2 port map ( Y=>nx30321, A0=>nx30325, A1=>
      max_calc_comparator_third_inp1_13);
   ix30340 : or03 port map ( Y=>nx30339, A0=>nx30122, A1=>nx36197, A2=>
      nx36069);
   ix30346 : or03 port map ( Y=>nx30345, A0=>nx30311, A1=>nx36197, A2=>
      nx36069);
   ix12221 : xnor2 port map ( Y=>nx12220, A0=>nx30336, A1=>nx30343);
   ix30350 : xnor2 port map ( Y=>nx30349, A0=>nx30353, A1=>
      max_calc_comparator_third_inp1_11);
   ix30368 : or03 port map ( Y=>nx30367, A0=>nx30107, A1=>nx36197, A2=>
      nx36069);
   ix30374 : or03 port map ( Y=>nx30373, A0=>nx30296, A1=>nx36197, A2=>
      nx36069);
   ix12265 : xnor2 port map ( Y=>nx12264, A0=>nx30364, A1=>nx30371);
   ix30378 : xnor2 port map ( Y=>nx30377, A0=>nx30381, A1=>
      max_calc_comparator_third_inp1_9);
   ix30396 : or03 port map ( Y=>nx30395, A0=>nx30092, A1=>nx36197, A2=>
      nx36069);
   ix30402 : or03 port map ( Y=>nx30401, A0=>nx30281, A1=>nx36197, A2=>
      nx35365);
   ix12309 : xnor2 port map ( Y=>nx12308, A0=>nx30392, A1=>nx30399);
   ix30406 : xnor2 port map ( Y=>nx30405, A0=>nx30409, A1=>
      max_calc_comparator_third_inp1_7);
   ix30424 : or03 port map ( Y=>nx30423, A0=>nx30077, A1=>nx36197, A2=>
      nx35365);
   ix30430 : or03 port map ( Y=>nx30429, A0=>nx30266, A1=>nx36199, A2=>
      nx35365);
   ix12353 : xnor2 port map ( Y=>nx12352, A0=>nx30420, A1=>nx30427);
   ix30434 : xnor2 port map ( Y=>nx30433, A0=>nx30437, A1=>
      max_calc_comparator_third_inp1_5);
   ix30452 : or03 port map ( Y=>nx30451, A0=>nx30062, A1=>nx36199, A2=>
      nx35365);
   ix30458 : or03 port map ( Y=>nx30457, A0=>nx30251, A1=>nx36199, A2=>
      nx35365);
   ix12397 : xnor2 port map ( Y=>nx12396, A0=>nx30448, A1=>nx30455);
   ix30462 : xnor2 port map ( Y=>nx30461, A0=>nx30465, A1=>
      max_calc_comparator_third_inp1_3);
   ix30480 : or03 port map ( Y=>nx30479, A0=>nx30047, A1=>nx36199, A2=>
      nx35365);
   ix30486 : or03 port map ( Y=>nx30485, A0=>nx30236, A1=>nx36199, A2=>
      nx36073);
   ix12441 : xnor2 port map ( Y=>nx12440, A0=>nx30476, A1=>nx30483);
   ix12463 : xnor2 port map ( Y=>nx12462, A0=>nx30491, A1=>nx30495);
   ix12689 : xnor2 port map ( Y=>nx12688, A0=>nx30506, A1=>nx30524);
   ix21614 : mux21_ni port map ( Y=>nx21613, A0=>label_6_output(15), A1=>
      label_6_input_15, S0=>nx36257);
   ix12625 : mux21_ni port map ( Y=>nx12624, A0=>nx12620, A1=>
      label_6_input_state_machine_15, S0=>nx35935);
   ix21604 : mux21_ni port map ( Y=>nx21603, A0=>
      label_6_input_state_machine_15, A1=>mdr_data_out(95), S0=>nx36219);
   ix30520 : xor2 port map ( Y=>nx30519, A0=>nx29921, A1=>label_6_output(15)
   );
   ix21644 : mux21_ni port map ( Y=>nx21643, A0=>label_5_output(15), A1=>
      label_5_input_15, S0=>nx36257);
   ix12667 : mux21_ni port map ( Y=>nx12666, A0=>nx12662, A1=>
      label_5_input_state_machine_15, S0=>nx35935);
   ix21634 : mux21_ni port map ( Y=>nx21633, A0=>
      label_5_input_state_machine_15, A1=>mdr_data_out(79), S0=>nx36219);
   ix30538 : xor2 port map ( Y=>nx30537, A0=>nx29480, A1=>label_5_output(15)
   );
   ix9537 : nand02 port map ( Y=>nx34913, A0=>nx36291, A1=>nx35869);
   ix9533 : nand04 port map ( Y=>nx34905, A0=>nx36291, A1=>nx35737, A2=>
      nx26203, A3=>nx35641);
   ix16897 : mux21_ni port map ( Y=>nx16896, A0=>max_calc_ans4_0, A1=>
      label_4_output(0), S0=>nx35979);
   ix14674 : mux21_ni port map ( Y=>nx14673, A0=>label_4_output(0), A1=>
      label_4_input_0, S0=>nx36257);
   ix14664 : mux21_ni port map ( Y=>nx14663, A0=>
      label_4_input_state_machine_0, A1=>mdr_data_out(48), S0=>nx36219);
   ix14654 : mux21_ni port map ( Y=>nx14653, A0=>nx35719, A1=>nx1722, S0=>
      nx35505);
   ix1723 : mux21_ni port map ( Y=>nx1722, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_3_1, S0=>nx36155);
   ix14644 : mux21_ni port map ( Y=>nx14643, A0=>
      booth_booth_integration_output_3_1, A1=>nx1710, S0=>nx35505);
   ix1711 : mux21_ni port map ( Y=>nx1710, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_3_2, S0=>nx36155);
   ix14634 : mux21_ni port map ( Y=>nx14633, A0=>
      booth_booth_integration_output_3_2, A1=>nx1698, S0=>nx35505);
   ix1699 : mux21_ni port map ( Y=>nx1698, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_3_3, S0=>nx36155);
   ix14624 : mux21_ni port map ( Y=>nx14623, A0=>
      booth_booth_integration_output_3_3, A1=>nx1686, S0=>nx35505);
   ix1687 : mux21_ni port map ( Y=>nx1686, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_3_4, S0=>nx36155);
   ix14614 : mux21_ni port map ( Y=>nx14613, A0=>
      booth_booth_integration_output_3_4, A1=>nx1674, S0=>nx35505);
   ix1675 : mux21_ni port map ( Y=>nx1674, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_3_5, S0=>nx36155);
   ix14604 : mux21_ni port map ( Y=>nx14603, A0=>
      booth_booth_integration_output_3_5, A1=>nx1662, S0=>nx35505);
   ix1663 : mux21_ni port map ( Y=>nx1662, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_3_6, S0=>nx36157);
   ix14594 : mux21_ni port map ( Y=>nx14593, A0=>
      booth_booth_integration_output_3_6, A1=>nx1650, S0=>nx35505);
   ix1651 : mux21_ni port map ( Y=>nx1650, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_3_7, S0=>nx36157);
   ix14584 : mux21_ni port map ( Y=>nx14583, A0=>
      booth_booth_integration_output_3_7, A1=>nx1638, S0=>nx36147);
   ix1639 : mux21_ni port map ( Y=>nx1638, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_3_8, S0=>nx36157);
   ix14574 : mux21_ni port map ( Y=>nx14573, A0=>
      booth_booth_integration_output_3_8, A1=>nx1626, S0=>nx36147);
   ix1627 : mux21_ni port map ( Y=>nx1626, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_3_9, S0=>nx36157);
   ix14564 : mux21_ni port map ( Y=>nx14563, A0=>
      booth_booth_integration_output_3_9, A1=>nx1614, S0=>nx36147);
   ix1615 : mux21_ni port map ( Y=>nx1614, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_3_10, S0=>nx36157);
   ix14554 : mux21_ni port map ( Y=>nx14553, A0=>
      booth_booth_integration_output_3_10, A1=>nx1602, S0=>nx36149);
   ix1603 : mux21_ni port map ( Y=>nx1602, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_3_11, S0=>nx36157);
   ix14544 : mux21_ni port map ( Y=>nx14543, A0=>
      booth_booth_integration_output_3_11, A1=>nx1590, S0=>nx36149);
   ix1591 : mux21_ni port map ( Y=>nx1590, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_3_12, S0=>nx36157);
   ix14534 : mux21_ni port map ( Y=>nx14533, A0=>
      booth_booth_integration_output_3_12, A1=>nx1578, S0=>nx36149);
   ix1579 : mux21_ni port map ( Y=>nx1578, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_3_13, S0=>nx36159);
   ix14524 : mux21_ni port map ( Y=>nx14523, A0=>
      booth_booth_integration_output_3_13, A1=>nx1566, S0=>nx36149);
   ix1567 : mux21_ni port map ( Y=>nx1566, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_3_14, S0=>nx36159);
   ix14514 : mux21_ni port map ( Y=>nx14513, A0=>
      booth_booth_integration_output_3_14, A1=>nx1554, S0=>nx36149);
   ix1555 : mux21_ni port map ( Y=>nx1554, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_3_15, S0=>nx36159);
   ix14504 : mux21 port map ( Y=>nx14503, A0=>nx30966, A1=>nx30608, S0=>
      nx36149);
   ix14154 : mux21_ni port map ( Y=>nx14153, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_0, A1=>nx34571, S0=>nx35831
   );
   ix14140 : and02 port map ( Y=>nx14139, A0=>nx36315, A1=>
      booth_booth_integrtaion_3_shift_Reg_count_0);
   ix14334 : mux21_ni port map ( Y=>nx14333, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_9, A1=>nx34557, S0=>nx35831
   );
   ix14324 : mux21_ni port map ( Y=>nx14323, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_8, S0=>nx36149);
   ix14314 : mux21_ni port map ( Y=>nx14313, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_8, S0=>nx35831);
   ix14304 : mux21_ni port map ( Y=>nx14303, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_7, S0=>nx36151);
   ix14294 : mux21_ni port map ( Y=>nx14293, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_7, S0=>nx35831);
   ix14284 : mux21_ni port map ( Y=>nx14283, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_6, S0=>nx36151);
   ix14274 : mux21_ni port map ( Y=>nx14273, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_6, S0=>nx35831);
   ix14264 : mux21_ni port map ( Y=>nx14263, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_5, S0=>nx36151);
   ix14254 : mux21_ni port map ( Y=>nx14253, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_5, S0=>nx35831);
   ix14244 : mux21_ni port map ( Y=>nx14243, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_4, S0=>nx36151);
   ix14234 : mux21_ni port map ( Y=>nx14233, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_4, S0=>nx35833);
   ix14224 : mux21_ni port map ( Y=>nx14223, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_3, S0=>nx36151);
   ix14214 : mux21_ni port map ( Y=>nx14213, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_3, S0=>nx35833);
   ix14204 : mux21_ni port map ( Y=>nx14203, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_2, S0=>nx36151);
   ix14194 : mux21_ni port map ( Y=>nx14193, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_2, S0=>nx35833);
   ix14184 : mux21_ni port map ( Y=>nx14183, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_1, S0=>nx36151);
   ix14174 : mux21_ni port map ( Y=>nx14173, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_3_shift_Reg_output_1, S0=>nx35833);
   ix14164 : mux21_ni port map ( Y=>nx14163, A0=>
      booth_booth_integrtaion_3_shift_Reg_count_1, A1=>nx34571, S0=>nx36153
   );
   ix995 : and02 port map ( Y=>nx994, A0=>nx30681, A1=>nx35719);
   ix30684 : or03 port map ( Y=>nx30683, A0=>nx30685, A1=>
      booth_booth_integrtaion_3_shift_reg_output_0, A2=>nx36315);
   ix14494 : mux21_ni port map ( Y=>nx14493, A0=>
      booth_booth_integrtaion_3_booth_output_16, A1=>nx1524, S0=>nx36153);
   ix1525 : nor02ii port map ( Y=>nx1524, A0=>nx30692, A1=>nx36159);
   ix1001 : nor02ii port map ( Y=>nx1000, A0=>nx30676, A1=>
      booth_booth_integrtaion_3_booth_output_16);
   ix1519 : xor2 port map ( Y=>nx12913, A0=>nx30698, A1=>nx30962);
   ix1507 : xor2 port map ( Y=>nx12915, A0=>nx30723, A1=>nx35511);
   ix14474 : mux21_ni port map ( Y=>nx14473, A0=>
      booth_booth_integrtaion_3_booth_output_18, A1=>nx1500, S0=>nx36153);
   ix1501 : nor02ii port map ( Y=>nx1500, A0=>nx30713, A1=>nx36159);
   ix1495 : xor2 port map ( Y=>nx12917, A0=>nx30728, A1=>nx30959);
   ix30745 : or02 port map ( Y=>nx30744, A0=>nx30681, A1=>nx35721);
   ix1483 : xor2 port map ( Y=>nx12919, A0=>nx30762, A1=>nx35513);
   ix14454 : mux21_ni port map ( Y=>nx14453, A0=>
      booth_booth_integrtaion_3_booth_output_20, A1=>nx1476, S0=>nx36153);
   ix1477 : nor02ii port map ( Y=>nx1476, A0=>nx30750, A1=>nx36159);
   ix1471 : xor2 port map ( Y=>nx12921, A0=>nx30767, A1=>nx30956);
   ix1459 : xor2 port map ( Y=>nx12922, A0=>nx30797, A1=>nx35515);
   ix14434 : mux21_ni port map ( Y=>nx14433, A0=>
      booth_booth_integrtaion_3_booth_output_22, A1=>nx1452, S0=>nx36153);
   ix1453 : nor02ii port map ( Y=>nx1452, A0=>nx30785, A1=>nx36159);
   ix1447 : xor2 port map ( Y=>nx12923, A0=>nx30802, A1=>nx30953);
   ix1435 : xor2 port map ( Y=>nx12925, A0=>nx30832, A1=>nx35517);
   ix14414 : mux21_ni port map ( Y=>nx14413, A0=>
      booth_booth_integrtaion_3_booth_output_24, A1=>nx1428, S0=>nx36153);
   ix1429 : nor02ii port map ( Y=>nx1428, A0=>nx30820, A1=>nx36161);
   ix1423 : xor2 port map ( Y=>nx12927, A0=>nx30837, A1=>nx30950);
   ix1411 : xor2 port map ( Y=>nx12929, A0=>nx30867, A1=>nx35519);
   ix14394 : mux21_ni port map ( Y=>nx14393, A0=>
      booth_booth_integrtaion_3_booth_output_26, A1=>nx1404, S0=>nx36153);
   ix1405 : nor02ii port map ( Y=>nx1404, A0=>nx30855, A1=>nx36161);
   ix1399 : xor2 port map ( Y=>nx12930, A0=>nx30872, A1=>nx30947);
   ix1387 : xor2 port map ( Y=>nx12931, A0=>nx30902, A1=>nx35521);
   ix14374 : mux21_ni port map ( Y=>nx14373, A0=>
      booth_booth_integrtaion_3_booth_output_28, A1=>nx1380, S0=>nx35503);
   ix1381 : nor02ii port map ( Y=>nx1380, A0=>nx30890, A1=>nx36161);
   ix1375 : xor2 port map ( Y=>nx12933, A0=>nx30907, A1=>nx30944);
   ix1363 : xor2 port map ( Y=>nx12935, A0=>nx30937, A1=>nx35523);
   ix14354 : mux21_ni port map ( Y=>nx14353, A0=>
      booth_booth_integrtaion_3_booth_output_31, A1=>nx1356, S0=>nx35503);
   ix1357 : nor02ii port map ( Y=>nx1356, A0=>nx30925, A1=>nx36161);
   ix1351 : xor2 port map ( Y=>nx1350, A0=>nx30937, A1=>nx30940);
   ix1537 : nor02ii port map ( Y=>nx1536, A0=>nx1000, A1=>nx36161);
   ix24244 : ao32 port map ( Y=>nx24243, A0=>nx35961, A1=>nx35647, A2=>
      nx36291, B0=>max_calc_ans4_0, B1=>nx35877);
   ix30987 : mux21 port map ( Y=>nx35647, A0=>nx31429, A1=>nx30990, S0=>
      nx35893);
   ix22234 : mux21_ni port map ( Y=>nx22233, A0=>label_7_output(0), A1=>
      label_7_input_0, S0=>nx36257);
   ix22224 : mux21_ni port map ( Y=>nx22223, A0=>
      label_7_input_state_machine_0, A1=>mdr_data_out(96), S0=>nx36219);
   ix22214 : mux21_ni port map ( Y=>nx22213, A0=>nx35771, A1=>nx13564, S0=>
      nx35531);
   ix13565 : mux21_ni port map ( Y=>nx13564, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_6_1, S0=>nx36171);
   ix22204 : mux21_ni port map ( Y=>nx22203, A0=>
      booth_booth_integration_output_6_1, A1=>nx13552, S0=>nx35531);
   ix13553 : mux21_ni port map ( Y=>nx13552, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_6_2, S0=>nx36171);
   ix22194 : mux21_ni port map ( Y=>nx22193, A0=>
      booth_booth_integration_output_6_2, A1=>nx13540, S0=>nx35531);
   ix13541 : mux21_ni port map ( Y=>nx13540, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_6_3, S0=>nx36171);
   ix22184 : mux21_ni port map ( Y=>nx22183, A0=>
      booth_booth_integration_output_6_3, A1=>nx13528, S0=>nx35531);
   ix13529 : mux21_ni port map ( Y=>nx13528, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_6_4, S0=>nx36171);
   ix22174 : mux21_ni port map ( Y=>nx22173, A0=>
      booth_booth_integration_output_6_4, A1=>nx13516, S0=>nx35531);
   ix13517 : mux21_ni port map ( Y=>nx13516, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_6_5, S0=>nx36171);
   ix22164 : mux21_ni port map ( Y=>nx22163, A0=>
      booth_booth_integration_output_6_5, A1=>nx13504, S0=>nx35531);
   ix13505 : mux21_ni port map ( Y=>nx13504, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_6_6, S0=>nx36173);
   ix22154 : mux21_ni port map ( Y=>nx22153, A0=>
      booth_booth_integration_output_6_6, A1=>nx13492, S0=>nx35531);
   ix13493 : mux21_ni port map ( Y=>nx13492, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_6_7, S0=>nx36173);
   ix22144 : mux21_ni port map ( Y=>nx22143, A0=>
      booth_booth_integration_output_6_7, A1=>nx13480, S0=>nx36163);
   ix13481 : mux21_ni port map ( Y=>nx13480, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_6_8, S0=>nx36173);
   ix22134 : mux21_ni port map ( Y=>nx22133, A0=>
      booth_booth_integration_output_6_8, A1=>nx13468, S0=>nx36163);
   ix13469 : mux21_ni port map ( Y=>nx13468, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_6_9, S0=>nx36173);
   ix22124 : mux21_ni port map ( Y=>nx22123, A0=>
      booth_booth_integration_output_6_9, A1=>nx13456, S0=>nx36163);
   ix13457 : mux21_ni port map ( Y=>nx13456, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_6_10, S0=>nx36173);
   ix22114 : mux21_ni port map ( Y=>nx22113, A0=>
      booth_booth_integration_output_6_10, A1=>nx13444, S0=>nx36165);
   ix13445 : mux21_ni port map ( Y=>nx13444, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_6_11, S0=>nx36173);
   ix22104 : mux21_ni port map ( Y=>nx22103, A0=>
      booth_booth_integration_output_6_11, A1=>nx13432, S0=>nx36165);
   ix13433 : mux21_ni port map ( Y=>nx13432, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_6_12, S0=>nx36173);
   ix22094 : mux21_ni port map ( Y=>nx22093, A0=>
      booth_booth_integration_output_6_12, A1=>nx13420, S0=>nx36165);
   ix13421 : mux21_ni port map ( Y=>nx13420, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_6_13, S0=>nx36175);
   ix22084 : mux21_ni port map ( Y=>nx22083, A0=>
      booth_booth_integration_output_6_13, A1=>nx13408, S0=>nx36165);
   ix13409 : mux21_ni port map ( Y=>nx13408, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_6_14, S0=>nx36175);
   ix22074 : mux21_ni port map ( Y=>nx22073, A0=>
      booth_booth_integration_output_6_14, A1=>nx13396, S0=>nx36165);
   ix13397 : mux21_ni port map ( Y=>nx13396, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_6_15, S0=>nx36175);
   ix22064 : mux21 port map ( Y=>nx22063, A0=>nx31409, A1=>nx31051, S0=>
      nx36165);
   ix21714 : mux21_ni port map ( Y=>nx21713, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_0, A1=>nx35011, S0=>nx35835
   );
   ix21700 : and02 port map ( Y=>nx21699, A0=>nx36357, A1=>
      booth_booth_integrtaion_6_shift_Reg_count_0);
   ix21894 : mux21_ni port map ( Y=>nx21893, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_9, A1=>nx34997, S0=>nx35835
   );
   ix21884 : mux21_ni port map ( Y=>nx21883, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_8, S0=>nx36165);
   ix21874 : mux21_ni port map ( Y=>nx21873, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_8, S0=>nx35835);
   ix21864 : mux21_ni port map ( Y=>nx21863, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_7, S0=>nx36167);
   ix21854 : mux21_ni port map ( Y=>nx21853, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_7, S0=>nx35835);
   ix21844 : mux21_ni port map ( Y=>nx21843, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_6, S0=>nx36167);
   ix21834 : mux21_ni port map ( Y=>nx21833, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_6, S0=>nx35835);
   ix21824 : mux21_ni port map ( Y=>nx21823, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_5, S0=>nx36167);
   ix21814 : mux21_ni port map ( Y=>nx21813, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_5, S0=>nx35835);
   ix21804 : mux21_ni port map ( Y=>nx21803, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_4, S0=>nx36167);
   ix21794 : mux21_ni port map ( Y=>nx21793, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_4, S0=>nx35837);
   ix21784 : mux21_ni port map ( Y=>nx21783, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_3, S0=>nx36167);
   ix21774 : mux21_ni port map ( Y=>nx21773, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_3, S0=>nx35837);
   ix21764 : mux21_ni port map ( Y=>nx21763, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_2, S0=>nx36167);
   ix21754 : mux21_ni port map ( Y=>nx21753, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_2, S0=>nx35837);
   ix21744 : mux21_ni port map ( Y=>nx21743, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_1, S0=>nx36167);
   ix21734 : mux21_ni port map ( Y=>nx21733, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_6_shift_Reg_output_1, S0=>nx35837);
   ix21724 : mux21_ni port map ( Y=>nx21723, A0=>
      booth_booth_integrtaion_6_shift_Reg_count_1, A1=>nx35011, S0=>nx36169
   );
   ix12837 : and02 port map ( Y=>nx12836, A0=>nx31124, A1=>nx35771);
   ix31127 : or03 port map ( Y=>nx31126, A0=>nx31128, A1=>
      booth_booth_integrtaion_6_shift_reg_output_0, A2=>nx36357);
   ix22054 : mux21_ni port map ( Y=>nx22053, A0=>
      booth_booth_integrtaion_6_booth_output_16, A1=>nx13366, S0=>nx36169);
   ix13367 : nor02ii port map ( Y=>nx13366, A0=>nx31135, A1=>nx36175);
   ix12843 : nor02ii port map ( Y=>nx12842, A0=>nx31119, A1=>
      booth_booth_integrtaion_6_booth_output_16);
   ix13361 : xor2 port map ( Y=>nx13296, A0=>nx31141, A1=>nx31405);
   ix13349 : xor2 port map ( Y=>nx13297, A0=>nx31166, A1=>nx35537);
   ix22034 : mux21_ni port map ( Y=>nx22033, A0=>
      booth_booth_integrtaion_6_booth_output_18, A1=>nx13342, S0=>nx36169);
   ix13343 : nor02ii port map ( Y=>nx13342, A0=>nx31156, A1=>nx36175);
   ix13337 : xor2 port map ( Y=>nx13298, A0=>nx31171, A1=>nx31402);
   ix31188 : or02 port map ( Y=>nx31187, A0=>nx31124, A1=>nx35773);
   ix13325 : xor2 port map ( Y=>nx13299, A0=>nx31205, A1=>nx35539);
   ix22014 : mux21_ni port map ( Y=>nx22013, A0=>
      booth_booth_integrtaion_6_booth_output_20, A1=>nx13318, S0=>nx36169);
   ix13319 : nor02ii port map ( Y=>nx13318, A0=>nx31193, A1=>nx36175);
   ix13313 : xor2 port map ( Y=>nx13300, A0=>nx31210, A1=>nx31399);
   ix13301 : xor2 port map ( Y=>nx13301, A0=>nx31240, A1=>nx35541);
   ix21994 : mux21_ni port map ( Y=>nx21993, A0=>
      booth_booth_integrtaion_6_booth_output_22, A1=>nx13294, S0=>nx36169);
   ix13295 : nor02ii port map ( Y=>nx13294, A0=>nx31228, A1=>nx36175);
   ix13289 : xor2 port map ( Y=>nx13303, A0=>nx31245, A1=>nx31396);
   ix13277 : xor2 port map ( Y=>nx13305, A0=>nx31275, A1=>nx35543);
   ix21974 : mux21_ni port map ( Y=>nx21973, A0=>
      booth_booth_integrtaion_6_booth_output_24, A1=>nx13270, S0=>nx36169);
   ix13271 : nor02ii port map ( Y=>nx13270, A0=>nx31263, A1=>nx36177);
   ix13265 : xor2 port map ( Y=>nx13307, A0=>nx31280, A1=>nx31393);
   ix13253 : xor2 port map ( Y=>nx13308, A0=>nx31310, A1=>nx35545);
   ix21954 : mux21_ni port map ( Y=>nx21953, A0=>
      booth_booth_integrtaion_6_booth_output_26, A1=>nx13246, S0=>nx36169);
   ix13247 : nor02ii port map ( Y=>nx13246, A0=>nx31298, A1=>nx36177);
   ix13241 : xor2 port map ( Y=>nx13309, A0=>nx31315, A1=>nx31390);
   ix13229 : xor2 port map ( Y=>nx13310, A0=>nx31345, A1=>nx35547);
   ix21934 : mux21_ni port map ( Y=>nx21933, A0=>
      booth_booth_integrtaion_6_booth_output_28, A1=>nx13222, S0=>nx35529);
   ix13223 : nor02ii port map ( Y=>nx13222, A0=>nx31333, A1=>nx36177);
   ix13217 : xor2 port map ( Y=>nx13311, A0=>nx31350, A1=>nx31387);
   ix13205 : xor2 port map ( Y=>nx13312, A0=>nx31380, A1=>nx35549);
   ix21914 : mux21_ni port map ( Y=>nx21913, A0=>
      booth_booth_integrtaion_6_booth_output_31, A1=>nx13198, S0=>nx35529);
   ix13199 : nor02ii port map ( Y=>nx13198, A0=>nx31368, A1=>nx36177);
   ix13193 : xor2 port map ( Y=>nx13192, A0=>nx31380, A1=>nx31383);
   ix13379 : nor02ii port map ( Y=>nx13378, A0=>nx12842, A1=>nx36177);
   ix23074 : mux21_ni port map ( Y=>nx23073, A0=>label_8_output(0), A1=>
      label_8_input_0, S0=>nx36257);
   ix23064 : mux21_ni port map ( Y=>nx23063, A0=>
      label_8_input_state_machine_0, A1=>mdr_data_out(112), S0=>nx36221);
   ix23054 : mux21_ni port map ( Y=>nx23053, A0=>nx35775, A1=>nx14880, S0=>
      nx35557);
   ix14881 : mux21_ni port map ( Y=>nx14880, A0=>mdr_data_out(0), A1=>
      booth_booth_integration_output_7_1, S0=>nx36187);
   ix23044 : mux21_ni port map ( Y=>nx23043, A0=>
      booth_booth_integration_output_7_1, A1=>nx14868, S0=>nx35557);
   ix14869 : mux21_ni port map ( Y=>nx14868, A0=>mdr_data_out(1), A1=>
      booth_booth_integration_output_7_2, S0=>nx36187);
   ix23034 : mux21_ni port map ( Y=>nx23033, A0=>
      booth_booth_integration_output_7_2, A1=>nx14856, S0=>nx35557);
   ix14857 : mux21_ni port map ( Y=>nx14856, A0=>mdr_data_out(2), A1=>
      booth_booth_integration_output_7_3, S0=>nx36187);
   ix23024 : mux21_ni port map ( Y=>nx23023, A0=>
      booth_booth_integration_output_7_3, A1=>nx14844, S0=>nx35557);
   ix14845 : mux21_ni port map ( Y=>nx14844, A0=>mdr_data_out(3), A1=>
      booth_booth_integration_output_7_4, S0=>nx36187);
   ix23014 : mux21_ni port map ( Y=>nx23013, A0=>
      booth_booth_integration_output_7_4, A1=>nx14832, S0=>nx35557);
   ix14833 : mux21_ni port map ( Y=>nx14832, A0=>mdr_data_out(4), A1=>
      booth_booth_integration_output_7_5, S0=>nx36187);
   ix23004 : mux21_ni port map ( Y=>nx23003, A0=>
      booth_booth_integration_output_7_5, A1=>nx14820, S0=>nx35557);
   ix14821 : mux21_ni port map ( Y=>nx14820, A0=>mdr_data_out(5), A1=>
      booth_booth_integration_output_7_6, S0=>nx36189);
   ix22994 : mux21_ni port map ( Y=>nx22993, A0=>
      booth_booth_integration_output_7_6, A1=>nx14808, S0=>nx35557);
   ix14809 : mux21_ni port map ( Y=>nx14808, A0=>mdr_data_out(6), A1=>
      booth_booth_integration_output_7_7, S0=>nx36189);
   ix22984 : mux21_ni port map ( Y=>nx22983, A0=>
      booth_booth_integration_output_7_7, A1=>nx14796, S0=>nx36179);
   ix14797 : mux21_ni port map ( Y=>nx14796, A0=>mdr_data_out(7), A1=>
      booth_booth_integration_output_7_8, S0=>nx36189);
   ix22974 : mux21_ni port map ( Y=>nx22973, A0=>
      booth_booth_integration_output_7_8, A1=>nx14784, S0=>nx36179);
   ix14785 : mux21_ni port map ( Y=>nx14784, A0=>mdr_data_out(8), A1=>
      booth_booth_integration_output_7_9, S0=>nx36189);
   ix22964 : mux21_ni port map ( Y=>nx22963, A0=>
      booth_booth_integration_output_7_9, A1=>nx14772, S0=>nx36179);
   ix14773 : mux21_ni port map ( Y=>nx14772, A0=>mdr_data_out(9), A1=>
      booth_booth_integration_output_7_10, S0=>nx36189);
   ix22954 : mux21_ni port map ( Y=>nx22953, A0=>
      booth_booth_integration_output_7_10, A1=>nx14760, S0=>nx36181);
   ix14761 : mux21_ni port map ( Y=>nx14760, A0=>mdr_data_out(10), A1=>
      booth_booth_integration_output_7_11, S0=>nx36189);
   ix22944 : mux21_ni port map ( Y=>nx22943, A0=>
      booth_booth_integration_output_7_11, A1=>nx14748, S0=>nx36181);
   ix14749 : mux21_ni port map ( Y=>nx14748, A0=>mdr_data_out(11), A1=>
      booth_booth_integration_output_7_12, S0=>nx36189);
   ix22934 : mux21_ni port map ( Y=>nx22933, A0=>
      booth_booth_integration_output_7_12, A1=>nx14736, S0=>nx36181);
   ix14737 : mux21_ni port map ( Y=>nx14736, A0=>mdr_data_out(12), A1=>
      booth_booth_integration_output_7_13, S0=>nx36191);
   ix22924 : mux21_ni port map ( Y=>nx22923, A0=>
      booth_booth_integration_output_7_13, A1=>nx14724, S0=>nx36181);
   ix14725 : mux21_ni port map ( Y=>nx14724, A0=>mdr_data_out(13), A1=>
      booth_booth_integration_output_7_14, S0=>nx36191);
   ix22914 : mux21_ni port map ( Y=>nx22913, A0=>
      booth_booth_integration_output_7_14, A1=>nx14712, S0=>nx36181);
   ix14713 : mux21_ni port map ( Y=>nx14712, A0=>mdr_data_out(14), A1=>
      booth_booth_integration_output_7_15, S0=>nx36191);
   ix22904 : mux21 port map ( Y=>nx22903, A0=>nx31848, A1=>nx31490, S0=>
      nx36181);
   ix22554 : mux21_ni port map ( Y=>nx22553, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_0, A1=>nx35043, S0=>nx35839
   );
   ix22540 : and02 port map ( Y=>nx22539, A0=>nx36361, A1=>
      booth_booth_integrtaion_7_shift_Reg_count_0);
   ix22734 : mux21_ni port map ( Y=>nx22733, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_9, A1=>nx35029, S0=>nx35839
   );
   ix22724 : mux21_ni port map ( Y=>nx22723, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_9, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_8, S0=>nx36181);
   ix22714 : mux21_ni port map ( Y=>nx22713, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_8, S0=>nx35839);
   ix22704 : mux21_ni port map ( Y=>nx22703, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_8, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_7, S0=>nx36183);
   ix22694 : mux21_ni port map ( Y=>nx22693, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_7, S0=>nx35839);
   ix22684 : mux21_ni port map ( Y=>nx22683, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_7, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_6, S0=>nx36183);
   ix22674 : mux21_ni port map ( Y=>nx22673, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_6, S0=>nx35839);
   ix22664 : mux21_ni port map ( Y=>nx22663, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_6, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_5, S0=>nx36183);
   ix22654 : mux21_ni port map ( Y=>nx22653, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_5, S0=>nx35839);
   ix22644 : mux21_ni port map ( Y=>nx22643, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_5, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_4, S0=>nx36183);
   ix22634 : mux21_ni port map ( Y=>nx22633, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_4, S0=>nx35841);
   ix22624 : mux21_ni port map ( Y=>nx22623, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_4, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_3, S0=>nx36183);
   ix22614 : mux21_ni port map ( Y=>nx22613, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_3, S0=>nx35841);
   ix22604 : mux21_ni port map ( Y=>nx22603, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_3, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_2, S0=>nx36183);
   ix22594 : mux21_ni port map ( Y=>nx22593, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_2, S0=>nx35841);
   ix22584 : mux21_ni port map ( Y=>nx22583, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_2, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_1, S0=>nx36183);
   ix22574 : mux21_ni port map ( Y=>nx22573, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_1, A1=>
      booth_booth_integrtaion_7_shift_Reg_output_1, S0=>nx35841);
   ix22564 : mux21_ni port map ( Y=>nx22563, A0=>
      booth_booth_integrtaion_7_shift_Reg_count_1, A1=>nx35043, S0=>nx36185
   );
   ix14153 : and02 port map ( Y=>nx14152, A0=>nx31563, A1=>nx35775);
   ix31566 : or03 port map ( Y=>nx31565, A0=>nx31567, A1=>
      booth_booth_integrtaion_7_shift_reg_output_0, A2=>nx36361);
   ix22894 : mux21_ni port map ( Y=>nx22893, A0=>
      booth_booth_integrtaion_7_booth_output_16, A1=>nx14682, S0=>nx36185);
   ix14683 : nor02ii port map ( Y=>nx14682, A0=>nx31574, A1=>nx36191);
   ix14159 : nor02ii port map ( Y=>nx14158, A0=>nx31558, A1=>
      booth_booth_integrtaion_7_booth_output_16);
   ix14677 : xor2 port map ( Y=>nx13334, A0=>nx31580, A1=>nx31844);
   ix14665 : xor2 port map ( Y=>nx13335, A0=>nx31605, A1=>nx35563);
   ix22874 : mux21_ni port map ( Y=>nx22873, A0=>
      booth_booth_integrtaion_7_booth_output_18, A1=>nx14658, S0=>nx36185);
   ix14659 : nor02ii port map ( Y=>nx14658, A0=>nx31595, A1=>nx36191);
   ix14653 : xor2 port map ( Y=>nx13336, A0=>nx31610, A1=>nx31841);
   ix31627 : or02 port map ( Y=>nx31626, A0=>nx31563, A1=>nx35777);
   ix14641 : xor2 port map ( Y=>nx13337, A0=>nx31644, A1=>nx35565);
   ix22854 : mux21_ni port map ( Y=>nx22853, A0=>
      booth_booth_integrtaion_7_booth_output_20, A1=>nx14634, S0=>nx36185);
   ix14635 : nor02ii port map ( Y=>nx14634, A0=>nx31632, A1=>nx36191);
   ix14629 : xor2 port map ( Y=>nx13339, A0=>nx31649, A1=>nx31838);
   ix14617 : xor2 port map ( Y=>nx13341, A0=>nx31679, A1=>nx35567);
   ix22834 : mux21_ni port map ( Y=>nx22833, A0=>
      booth_booth_integrtaion_7_booth_output_22, A1=>nx14610, S0=>nx36185);
   ix14611 : nor02ii port map ( Y=>nx14610, A0=>nx31667, A1=>nx36191);
   ix14605 : xor2 port map ( Y=>nx13343, A0=>nx31684, A1=>nx31835);
   ix14593 : xor2 port map ( Y=>nx13344, A0=>nx31714, A1=>nx35569);
   ix22814 : mux21_ni port map ( Y=>nx22813, A0=>
      booth_booth_integrtaion_7_booth_output_24, A1=>nx14586, S0=>nx36185);
   ix14587 : nor02ii port map ( Y=>nx14586, A0=>nx31702, A1=>nx36193);
   ix14581 : xor2 port map ( Y=>nx13345, A0=>nx31719, A1=>nx31832);
   ix14569 : xor2 port map ( Y=>nx13346, A0=>nx31749, A1=>nx35571);
   ix22794 : mux21_ni port map ( Y=>nx22793, A0=>
      booth_booth_integrtaion_7_booth_output_26, A1=>nx14562, S0=>nx36185);
   ix14563 : nor02ii port map ( Y=>nx14562, A0=>nx31737, A1=>nx36193);
   ix14557 : xor2 port map ( Y=>nx13347, A0=>nx31754, A1=>nx31829);
   ix14545 : xor2 port map ( Y=>nx13348, A0=>nx31784, A1=>nx35573);
   ix22774 : mux21_ni port map ( Y=>nx22773, A0=>
      booth_booth_integrtaion_7_booth_output_28, A1=>nx14538, S0=>nx35555);
   ix14539 : nor02ii port map ( Y=>nx14538, A0=>nx31772, A1=>nx36193);
   ix14533 : xor2 port map ( Y=>nx13349, A0=>nx31789, A1=>nx31826);
   ix14521 : xor2 port map ( Y=>nx13351, A0=>nx31819, A1=>nx35575);
   ix22754 : mux21_ni port map ( Y=>nx22753, A0=>
      booth_booth_integrtaion_7_booth_output_31, A1=>nx14514, S0=>nx35555);
   ix14515 : nor02ii port map ( Y=>nx14514, A0=>nx31807, A1=>nx36193);
   ix14509 : xor2 port map ( Y=>nx14508, A0=>nx31819, A1=>nx31822);
   ix14695 : nor02ii port map ( Y=>nx14694, A0=>nx14158, A1=>nx36193);
   ix31873 : or03 port map ( Y=>nx31872, A0=>nx32056, A1=>nx36199, A2=>
      nx36073);
   ix23344 : mux21_ni port map ( Y=>nx23343, A0=>label_8_output(14), A1=>
      label_8_input_14, S0=>nx36259);
   ix15339 : mux21_ni port map ( Y=>nx15338, A0=>nx15334, A1=>
      label_8_input_state_machine_14, S0=>nx35937);
   ix22524 : mux21_ni port map ( Y=>nx22523, A0=>
      label_8_input_state_machine_14, A1=>mdr_data_out(126), S0=>nx36221);
   ix23334 : mux21_ni port map ( Y=>nx23333, A0=>label_8_output(13), A1=>
      label_8_input_13, S0=>nx36259);
   ix15313 : mux21_ni port map ( Y=>nx15312, A0=>nx15308, A1=>
      label_8_input_state_machine_13, S0=>nx35937);
   ix23324 : mux21_ni port map ( Y=>nx23323, A0=>
      label_8_input_state_machine_13, A1=>mdr_data_out(125), S0=>nx36221);
   ix23294 : mux21_ni port map ( Y=>nx23293, A0=>label_8_output(11), A1=>
      label_8_input_11, S0=>nx36259);
   ix15249 : mux21_ni port map ( Y=>nx15248, A0=>nx15244, A1=>
      label_8_input_state_machine_11, S0=>nx35937);
   ix23284 : mux21_ni port map ( Y=>nx23283, A0=>
      label_8_input_state_machine_11, A1=>mdr_data_out(123), S0=>nx36221);
   ix23254 : mux21_ni port map ( Y=>nx23253, A0=>label_8_output(9), A1=>
      label_8_input_9, S0=>nx36259);
   ix15185 : mux21_ni port map ( Y=>nx15184, A0=>nx15180, A1=>
      label_8_input_state_machine_9, S0=>nx35937);
   ix23244 : mux21_ni port map ( Y=>nx23243, A0=>
      label_8_input_state_machine_9, A1=>mdr_data_out(121), S0=>nx36221);
   ix23214 : mux21_ni port map ( Y=>nx23213, A0=>label_8_output(7), A1=>
      label_8_input_7, S0=>nx36259);
   ix15121 : mux21_ni port map ( Y=>nx15120, A0=>nx15116, A1=>
      label_8_input_state_machine_7, S0=>nx35937);
   ix23204 : mux21_ni port map ( Y=>nx23203, A0=>
      label_8_input_state_machine_7, A1=>mdr_data_out(119), S0=>nx36221);
   ix23174 : mux21_ni port map ( Y=>nx23173, A0=>label_8_output(5), A1=>
      label_8_input_5, S0=>nx36259);
   ix15057 : mux21_ni port map ( Y=>nx15056, A0=>nx15052, A1=>
      label_8_input_state_machine_5, S0=>nx35937);
   ix23164 : mux21_ni port map ( Y=>nx23163, A0=>
      label_8_input_state_machine_5, A1=>mdr_data_out(117), S0=>nx36221);
   ix23134 : mux21_ni port map ( Y=>nx23133, A0=>label_8_output(3), A1=>
      label_8_input_3, S0=>nx36259);
   ix14993 : mux21_ni port map ( Y=>nx14992, A0=>nx14988, A1=>
      label_8_input_state_machine_3, S0=>nx35935);
   ix23124 : mux21_ni port map ( Y=>nx23123, A0=>
      label_8_input_state_machine_3, A1=>mdr_data_out(115), S0=>nx36223);
   ix23094 : mux21_ni port map ( Y=>nx23093, A0=>label_8_output(1), A1=>
      label_8_input_1, S0=>nx36261);
   ix14929 : mux21_ni port map ( Y=>nx14928, A0=>nx14924, A1=>
      label_8_input_state_machine_1, S0=>nx35935);
   ix23084 : mux21_ni port map ( Y=>nx23083, A0=>
      label_8_input_state_machine_1, A1=>mdr_data_out(113), S0=>nx36223);
   ix31965 : xnor2 port map ( Y=>nx31964, A0=>nx31862, A1=>nx31974);
   ix23114 : mux21_ni port map ( Y=>nx23113, A0=>label_8_output(2), A1=>
      label_8_input_2, S0=>nx36261);
   ix14961 : mux21_ni port map ( Y=>nx14960, A0=>nx14956, A1=>
      label_8_input_state_machine_2, S0=>nx35167);
   ix23104 : mux21_ni port map ( Y=>nx23103, A0=>
      label_8_input_state_machine_2, A1=>mdr_data_out(114), S0=>nx36223);
   ix31980 : xnor2 port map ( Y=>nx31979, A0=>nx31860, A1=>nx31989);
   ix23154 : mux21_ni port map ( Y=>nx23153, A0=>label_8_output(4), A1=>
      label_8_input_4, S0=>nx36261);
   ix15025 : mux21_ni port map ( Y=>nx15024, A0=>nx15020, A1=>
      label_8_input_state_machine_4, S0=>nx35167);
   ix23144 : mux21_ni port map ( Y=>nx23143, A0=>
      label_8_input_state_machine_4, A1=>mdr_data_out(116), S0=>nx36223);
   ix31995 : xnor2 port map ( Y=>nx31994, A0=>nx31858, A1=>nx32004);
   ix23194 : mux21_ni port map ( Y=>nx23193, A0=>label_8_output(6), A1=>
      label_8_input_6, S0=>nx36261);
   ix15089 : mux21_ni port map ( Y=>nx15088, A0=>nx15084, A1=>
      label_8_input_state_machine_6, S0=>nx35937);
   ix23184 : mux21_ni port map ( Y=>nx23183, A0=>
      label_8_input_state_machine_6, A1=>mdr_data_out(118), S0=>nx36223);
   ix32010 : xnor2 port map ( Y=>nx32009, A0=>nx31856, A1=>nx32019);
   ix23234 : mux21_ni port map ( Y=>nx23233, A0=>label_8_output(8), A1=>
      label_8_input_8, S0=>nx36261);
   ix15153 : mux21_ni port map ( Y=>nx15152, A0=>nx15148, A1=>
      label_8_input_state_machine_8, S0=>nx35939);
   ix23224 : mux21_ni port map ( Y=>nx23223, A0=>
      label_8_input_state_machine_8, A1=>mdr_data_out(120), S0=>nx36223);
   ix32025 : xnor2 port map ( Y=>nx32024, A0=>nx31854, A1=>nx32034);
   ix23274 : mux21_ni port map ( Y=>nx23273, A0=>label_8_output(10), A1=>
      label_8_input_10, S0=>nx36261);
   ix15217 : mux21_ni port map ( Y=>nx15216, A0=>nx15212, A1=>
      label_8_input_state_machine_10, S0=>nx35939);
   ix23264 : mux21_ni port map ( Y=>nx23263, A0=>
      label_8_input_state_machine_10, A1=>mdr_data_out(122), S0=>nx36223);
   ix32040 : xnor2 port map ( Y=>nx32039, A0=>nx31852, A1=>nx32049);
   ix23314 : mux21_ni port map ( Y=>nx23313, A0=>label_8_output(12), A1=>
      label_8_input_12, S0=>nx36261);
   ix15281 : mux21_ni port map ( Y=>nx15280, A0=>nx15276, A1=>
      label_8_input_state_machine_12, S0=>nx35939);
   ix23304 : mux21_ni port map ( Y=>nx23303, A0=>
      label_8_input_state_machine_12, A1=>mdr_data_out(124), S0=>nx35597);
   ix32055 : xnor2 port map ( Y=>nx32054, A0=>nx31850, A1=>nx32056);
   ix32062 : or03 port map ( Y=>nx32061, A0=>nx32245, A1=>nx36125, A2=>
      nx36073);
   ix22504 : mux21_ni port map ( Y=>nx22503, A0=>label_7_output(14), A1=>
      label_7_input_14, S0=>nx36263);
   ix14023 : mux21_ni port map ( Y=>nx14022, A0=>nx14018, A1=>
      label_7_input_state_machine_14, S0=>nx35939);
   ix21684 : mux21_ni port map ( Y=>nx21683, A0=>
      label_7_input_state_machine_14, A1=>mdr_data_out(110), S0=>nx35597);
   ix22494 : mux21_ni port map ( Y=>nx22493, A0=>label_7_output(13), A1=>
      label_7_input_13, S0=>nx36263);
   ix13997 : mux21_ni port map ( Y=>nx13996, A0=>nx13992, A1=>
      label_7_input_state_machine_13, S0=>nx35939);
   ix22484 : mux21_ni port map ( Y=>nx22483, A0=>
      label_7_input_state_machine_13, A1=>mdr_data_out(109), S0=>nx35597);
   ix22454 : mux21_ni port map ( Y=>nx22453, A0=>label_7_output(11), A1=>
      label_7_input_11, S0=>nx36263);
   ix13933 : mux21_ni port map ( Y=>nx13932, A0=>nx13928, A1=>
      label_7_input_state_machine_11, S0=>nx35939);
   ix22444 : mux21_ni port map ( Y=>nx22443, A0=>
      label_7_input_state_machine_11, A1=>mdr_data_out(107), S0=>nx35597);
   ix22414 : mux21_ni port map ( Y=>nx22413, A0=>label_7_output(9), A1=>
      label_7_input_9, S0=>nx36263);
   ix13869 : mux21_ni port map ( Y=>nx13868, A0=>nx13864, A1=>
      label_7_input_state_machine_9, S0=>nx35939);
   ix22404 : mux21_ni port map ( Y=>nx22403, A0=>
      label_7_input_state_machine_9, A1=>mdr_data_out(105), S0=>nx35597);
   ix22374 : mux21_ni port map ( Y=>nx22373, A0=>label_7_output(7), A1=>
      label_7_input_7, S0=>nx36263);
   ix13805 : mux21_ni port map ( Y=>nx13804, A0=>nx13800, A1=>
      label_7_input_state_machine_7, S0=>nx35941);
   ix22364 : mux21_ni port map ( Y=>nx22363, A0=>
      label_7_input_state_machine_7, A1=>mdr_data_out(103), S0=>nx35597);
   ix22334 : mux21_ni port map ( Y=>nx22333, A0=>label_7_output(5), A1=>
      label_7_input_5, S0=>nx36263);
   ix13741 : mux21_ni port map ( Y=>nx13740, A0=>nx13736, A1=>
      label_7_input_state_machine_5, S0=>nx35941);
   ix22324 : mux21_ni port map ( Y=>nx22323, A0=>
      label_7_input_state_machine_5, A1=>mdr_data_out(101), S0=>nx35597);
   ix22294 : mux21_ni port map ( Y=>nx22293, A0=>label_7_output(3), A1=>
      label_7_input_3, S0=>nx36263);
   ix13677 : mux21_ni port map ( Y=>nx13676, A0=>nx13672, A1=>
      label_7_input_state_machine_3, S0=>nx35941);
   ix22284 : mux21_ni port map ( Y=>nx22283, A0=>
      label_7_input_state_machine_3, A1=>mdr_data_out(99), S0=>nx36225);
   ix22254 : mux21_ni port map ( Y=>nx22253, A0=>label_7_output(1), A1=>
      label_7_input_1, S0=>nx35605);
   ix13613 : mux21_ni port map ( Y=>nx13612, A0=>nx13608, A1=>
      label_7_input_state_machine_1, S0=>nx35941);
   ix22244 : mux21_ni port map ( Y=>nx22243, A0=>
      label_7_input_state_machine_1, A1=>mdr_data_out(97), S0=>nx36225);
   ix32154 : xnor2 port map ( Y=>nx32153, A0=>nx31423, A1=>nx32163);
   ix22274 : mux21_ni port map ( Y=>nx22273, A0=>label_7_output(2), A1=>
      label_7_input_2, S0=>nx35605);
   ix13645 : mux21_ni port map ( Y=>nx13644, A0=>nx13640, A1=>
      label_7_input_state_machine_2, S0=>nx35941);
   ix22264 : mux21_ni port map ( Y=>nx22263, A0=>
      label_7_input_state_machine_2, A1=>mdr_data_out(98), S0=>nx36225);
   ix32169 : xnor2 port map ( Y=>nx32168, A0=>nx31421, A1=>nx32178);
   ix22314 : mux21_ni port map ( Y=>nx22313, A0=>label_7_output(4), A1=>
      label_7_input_4, S0=>nx35605);
   ix13709 : mux21_ni port map ( Y=>nx13708, A0=>nx13704, A1=>
      label_7_input_state_machine_4, S0=>nx35941);
   ix22304 : mux21_ni port map ( Y=>nx22303, A0=>
      label_7_input_state_machine_4, A1=>mdr_data_out(100), S0=>nx36225);
   ix32184 : xnor2 port map ( Y=>nx32183, A0=>nx31419, A1=>nx32193);
   ix22354 : mux21_ni port map ( Y=>nx22353, A0=>label_7_output(6), A1=>
      label_7_input_6, S0=>nx35605);
   ix13773 : mux21_ni port map ( Y=>nx13772, A0=>nx13768, A1=>
      label_7_input_state_machine_6, S0=>nx35941);
   ix22344 : mux21_ni port map ( Y=>nx22343, A0=>
      label_7_input_state_machine_6, A1=>mdr_data_out(102), S0=>nx36225);
   ix32199 : xnor2 port map ( Y=>nx32198, A0=>nx31417, A1=>nx32208);
   ix22394 : mux21_ni port map ( Y=>nx22393, A0=>label_7_output(8), A1=>
      label_7_input_8, S0=>nx35605);
   ix13837 : mux21_ni port map ( Y=>nx13836, A0=>nx13832, A1=>
      label_7_input_state_machine_8, S0=>nx35943);
   ix22384 : mux21_ni port map ( Y=>nx22383, A0=>
      label_7_input_state_machine_8, A1=>mdr_data_out(104), S0=>nx36225);
   ix32214 : xnor2 port map ( Y=>nx32213, A0=>nx31415, A1=>nx32223);
   ix22434 : mux21_ni port map ( Y=>nx22433, A0=>label_7_output(10), A1=>
      label_7_input_10, S0=>nx35605);
   ix13901 : mux21_ni port map ( Y=>nx13900, A0=>nx13896, A1=>
      label_7_input_state_machine_10, S0=>nx35943);
   ix22424 : mux21_ni port map ( Y=>nx22423, A0=>
      label_7_input_state_machine_10, A1=>mdr_data_out(106), S0=>nx36225);
   ix32229 : xnor2 port map ( Y=>nx32228, A0=>nx31413, A1=>nx32238);
   ix22474 : mux21_ni port map ( Y=>nx22473, A0=>label_7_output(12), A1=>
      label_7_input_12, S0=>nx35605);
   ix13965 : mux21_ni port map ( Y=>nx13964, A0=>nx13960, A1=>
      label_7_input_state_machine_12, S0=>nx35943);
   ix22464 : mux21_ni port map ( Y=>nx22463, A0=>
      label_7_input_state_machine_12, A1=>mdr_data_out(108), S0=>nx36227);
   ix32244 : xnor2 port map ( Y=>nx32243, A0=>nx31411, A1=>nx32245);
   ix15361 : xnor2 port map ( Y=>nx15360, A0=>nx31869, A1=>nx32059);
   ix32249 : xnor2 port map ( Y=>nx32248, A0=>nx32252, A1=>
      max_calc_comparator_fourth_inp1_13);
   ix32267 : or03 port map ( Y=>nx32266, A0=>nx32049, A1=>nx36125, A2=>
      nx36073);
   ix32273 : or03 port map ( Y=>nx32272, A0=>nx32238, A1=>nx36125, A2=>
      nx36073);
   ix15405 : xnor2 port map ( Y=>nx15404, A0=>nx32263, A1=>nx32270);
   ix32277 : xnor2 port map ( Y=>nx32276, A0=>nx32280, A1=>
      max_calc_comparator_fourth_inp1_11);
   ix32295 : or03 port map ( Y=>nx32294, A0=>nx32034, A1=>nx36127, A2=>
      nx36073);
   ix32301 : or03 port map ( Y=>nx32300, A0=>nx32223, A1=>nx36127, A2=>
      nx36073);
   ix15449 : xnor2 port map ( Y=>nx15448, A0=>nx32291, A1=>nx32298);
   ix32305 : xnor2 port map ( Y=>nx32304, A0=>nx32308, A1=>
      max_calc_comparator_fourth_inp1_9);
   ix32323 : or03 port map ( Y=>nx32322, A0=>nx32019, A1=>nx36127, A2=>
      nx35367);
   ix32329 : or03 port map ( Y=>nx32328, A0=>nx32208, A1=>nx36127, A2=>
      nx35367);
   ix15493 : xnor2 port map ( Y=>nx15492, A0=>nx32319, A1=>nx32326);
   ix32333 : xnor2 port map ( Y=>nx32332, A0=>nx32336, A1=>
      max_calc_comparator_fourth_inp1_7);
   ix32351 : or03 port map ( Y=>nx32350, A0=>nx32004, A1=>nx36127, A2=>
      nx35369);
   ix32357 : or03 port map ( Y=>nx32356, A0=>nx32193, A1=>nx36127, A2=>
      nx35369);
   ix15537 : xnor2 port map ( Y=>nx15536, A0=>nx32347, A1=>nx32354);
   ix32361 : xnor2 port map ( Y=>nx32360, A0=>nx32364, A1=>
      max_calc_comparator_fourth_inp1_5);
   ix32379 : or03 port map ( Y=>nx32378, A0=>nx31989, A1=>nx36127, A2=>
      nx35369);
   ix32385 : or03 port map ( Y=>nx32384, A0=>nx32178, A1=>nx36129, A2=>
      nx35369);
   ix15581 : xnor2 port map ( Y=>nx15580, A0=>nx32375, A1=>nx32382);
   ix32389 : xnor2 port map ( Y=>nx32388, A0=>nx32392, A1=>
      max_calc_comparator_fourth_inp1_3);
   ix32407 : or03 port map ( Y=>nx32406, A0=>nx31974, A1=>nx36129, A2=>
      nx35369);
   ix32413 : or03 port map ( Y=>nx32412, A0=>nx32163, A1=>nx36129, A2=>
      nx35369);
   ix15625 : xnor2 port map ( Y=>nx15624, A0=>nx32403, A1=>nx32410);
   ix15647 : xnor2 port map ( Y=>nx15646, A0=>nx32418, A1=>nx32422);
   ix15873 : xnor2 port map ( Y=>nx15872, A0=>nx32433, A1=>nx32451);
   ix23654 : mux21_ni port map ( Y=>nx23653, A0=>label_8_output(15), A1=>
      label_8_input_15, S0=>nx36265);
   ix15809 : mux21_ni port map ( Y=>nx15808, A0=>nx15804, A1=>
      label_8_input_state_machine_15, S0=>nx35943);
   ix23644 : mux21_ni port map ( Y=>nx23643, A0=>
      label_8_input_state_machine_15, A1=>mdr_data_out(127), S0=>nx36227);
   ix32447 : xor2 port map ( Y=>nx32446, A0=>nx31848, A1=>label_8_output(15)
   );
   ix32454 : or03 port map ( Y=>nx32453, A0=>nx35649, A1=>nx36129, A2=>
      nx35369);
   ix35648 : inv01 port map ( Y=>nx35649, A=>label_7_output(15));
   ix23684 : mux21_ni port map ( Y=>nx23683, A0=>label_7_output(15), A1=>
      label_7_input_15, S0=>nx36265);
   ix15851 : mux21_ni port map ( Y=>nx15850, A0=>nx15846, A1=>
      label_7_input_state_machine_15, S0=>nx35943);
   ix23674 : mux21_ni port map ( Y=>nx23673, A0=>
      label_7_input_state_machine_15, A1=>mdr_data_out(111), S0=>nx36227);
   ix32465 : xor2 port map ( Y=>nx32464, A0=>nx31409, A1=>label_7_output(15)
   );
   ix15897 : mux21 port map ( Y=>nx15896, A0=>nx32665, A1=>nx32660, S0=>
      nx35979);
   ix14954 : mux21_ni port map ( Y=>nx14953, A0=>label_4_output(14), A1=>
      label_4_input_14, S0=>nx36265);
   ix2187 : mux21_ni port map ( Y=>nx2186, A0=>nx2182, A1=>
      label_4_input_state_machine_14, S0=>nx35943);
   ix14944 : mux21_ni port map ( Y=>nx14943, A0=>
      label_4_input_state_machine_14, A1=>mdr_data_out(62), S0=>nx36227);
   ix14934 : mux21_ni port map ( Y=>nx14933, A0=>label_4_output(13), A1=>
      label_4_input_13, S0=>nx36265);
   ix2155 : mux21_ni port map ( Y=>nx2154, A0=>nx2150, A1=>
      label_4_input_state_machine_13, S0=>nx35943);
   ix14924 : mux21_ni port map ( Y=>nx14923, A0=>
      label_4_input_state_machine_13, A1=>mdr_data_out(61), S0=>nx36227);
   ix14894 : mux21_ni port map ( Y=>nx14893, A0=>label_4_output(11), A1=>
      label_4_input_11, S0=>nx36265);
   ix2091 : mux21_ni port map ( Y=>nx2090, A0=>nx2086, A1=>
      label_4_input_state_machine_11, S0=>nx35945);
   ix14884 : mux21_ni port map ( Y=>nx14883, A0=>
      label_4_input_state_machine_11, A1=>mdr_data_out(59), S0=>nx36227);
   ix14854 : mux21_ni port map ( Y=>nx14853, A0=>label_4_output(9), A1=>
      label_4_input_9, S0=>nx36265);
   ix2027 : mux21_ni port map ( Y=>nx2026, A0=>nx2022, A1=>
      label_4_input_state_machine_9, S0=>nx35945);
   ix14844 : mux21_ni port map ( Y=>nx14843, A0=>
      label_4_input_state_machine_9, A1=>mdr_data_out(57), S0=>nx36227);
   ix14814 : mux21_ni port map ( Y=>nx14813, A0=>label_4_output(7), A1=>
      label_4_input_7, S0=>nx36265);
   ix1963 : mux21_ni port map ( Y=>nx1962, A0=>nx1958, A1=>
      label_4_input_state_machine_7, S0=>nx35945);
   ix14804 : mux21_ni port map ( Y=>nx14803, A0=>
      label_4_input_state_machine_7, A1=>mdr_data_out(55), S0=>nx36229);
   ix14774 : mux21_ni port map ( Y=>nx14773, A0=>label_4_output(5), A1=>
      label_4_input_5, S0=>nx36267);
   ix1899 : mux21_ni port map ( Y=>nx1898, A0=>nx1894, A1=>
      label_4_input_state_machine_5, S0=>nx35945);
   ix14764 : mux21_ni port map ( Y=>nx14763, A0=>
      label_4_input_state_machine_5, A1=>mdr_data_out(53), S0=>nx36229);
   ix14734 : mux21_ni port map ( Y=>nx14733, A0=>label_4_output(3), A1=>
      label_4_input_3, S0=>nx36267);
   ix1835 : mux21_ni port map ( Y=>nx1834, A0=>nx1830, A1=>
      label_4_input_state_machine_3, S0=>nx35945);
   ix14724 : mux21_ni port map ( Y=>nx14723, A0=>
      label_4_input_state_machine_3, A1=>mdr_data_out(51), S0=>nx36229);
   ix14694 : mux21_ni port map ( Y=>nx14693, A0=>label_4_output(1), A1=>
      label_4_input_1, S0=>nx36267);
   ix1771 : mux21_ni port map ( Y=>nx1770, A0=>nx1766, A1=>
      label_4_input_state_machine_1, S0=>nx35945);
   ix14684 : mux21_ni port map ( Y=>nx14683, A0=>
      label_4_input_state_machine_1, A1=>mdr_data_out(49), S0=>nx36229);
   ix32569 : xnor2 port map ( Y=>nx32568, A0=>nx30980, A1=>nx32578);
   ix14714 : mux21_ni port map ( Y=>nx14713, A0=>label_4_output(2), A1=>
      label_4_input_2, S0=>nx36267);
   ix1803 : mux21_ni port map ( Y=>nx1802, A0=>nx1798, A1=>
      label_4_input_state_machine_2, S0=>nx35945);
   ix14704 : mux21_ni port map ( Y=>nx14703, A0=>
      label_4_input_state_machine_2, A1=>mdr_data_out(50), S0=>nx36229);
   ix32584 : xnor2 port map ( Y=>nx32583, A0=>nx30978, A1=>nx32593);
   ix14754 : mux21_ni port map ( Y=>nx14753, A0=>label_4_output(4), A1=>
      label_4_input_4, S0=>nx36267);
   ix1867 : mux21_ni port map ( Y=>nx1866, A0=>nx1862, A1=>
      label_4_input_state_machine_4, S0=>nx35947);
   ix14744 : mux21_ni port map ( Y=>nx14743, A0=>
      label_4_input_state_machine_4, A1=>mdr_data_out(52), S0=>nx36229);
   ix32599 : xnor2 port map ( Y=>nx32598, A0=>nx30976, A1=>nx32608);
   ix14794 : mux21_ni port map ( Y=>nx14793, A0=>label_4_output(6), A1=>
      label_4_input_6, S0=>nx36267);
   ix1931 : mux21_ni port map ( Y=>nx1930, A0=>nx1926, A1=>
      label_4_input_state_machine_6, S0=>nx35947);
   ix14784 : mux21_ni port map ( Y=>nx14783, A0=>
      label_4_input_state_machine_6, A1=>mdr_data_out(54), S0=>nx36229);
   ix32614 : xnor2 port map ( Y=>nx32613, A0=>nx30974, A1=>nx32623);
   ix14834 : mux21_ni port map ( Y=>nx14833, A0=>label_4_output(8), A1=>
      label_4_input_8, S0=>nx36267);
   ix1995 : mux21_ni port map ( Y=>nx1994, A0=>nx1990, A1=>
      label_4_input_state_machine_8, S0=>nx35947);
   ix14824 : mux21_ni port map ( Y=>nx14823, A0=>
      label_4_input_state_machine_8, A1=>mdr_data_out(56), S0=>nx36231);
   ix32629 : xnor2 port map ( Y=>nx32628, A0=>nx30972, A1=>nx32638);
   ix14874 : mux21_ni port map ( Y=>nx14873, A0=>label_4_output(10), A1=>
      label_4_input_10, S0=>nx36269);
   ix2059 : mux21_ni port map ( Y=>nx2058, A0=>nx2054, A1=>
      label_4_input_state_machine_10, S0=>nx35947);
   ix14864 : mux21_ni port map ( Y=>nx14863, A0=>
      label_4_input_state_machine_10, A1=>mdr_data_out(58), S0=>nx36231);
   ix32644 : xnor2 port map ( Y=>nx32643, A0=>nx30970, A1=>nx32653);
   ix14914 : mux21_ni port map ( Y=>nx14913, A0=>label_4_output(12), A1=>
      label_4_input_12, S0=>nx36269);
   ix2123 : mux21_ni port map ( Y=>nx2122, A0=>nx2118, A1=>
      label_4_input_state_machine_12, S0=>nx35947);
   ix14904 : mux21_ni port map ( Y=>nx14903, A0=>
      label_4_input_state_machine_12, A1=>mdr_data_out(60), S0=>nx36231);
   ix32659 : xnor2 port map ( Y=>nx32658, A0=>nx30968, A1=>nx32660);
   ix23704 : ao32 port map ( Y=>nx23703, A0=>nx35961, A1=>nx35651, A2=>
      nx36291, B0=>max_calc_ans4_14, B1=>nx35877);
   ix32664 : mux21 port map ( Y=>nx35651, A0=>nx31869, A1=>nx32059, S0=>
      nx35893);
   ix12713 : mux21 port map ( Y=>nx12712, A0=>nx32861, A1=>nx32856, S0=>
      nx35979);
   ix15804 : mux21_ni port map ( Y=>nx15803, A0=>label_3_output(14), A1=>
      label_3_input_14, S0=>nx36269);
   ix3525 : mux21_ni port map ( Y=>nx3524, A0=>nx3520, A1=>
      label_3_input_state_machine_14, S0=>nx35949);
   ix15794 : mux21_ni port map ( Y=>nx15793, A0=>
      label_3_input_state_machine_14, A1=>mdr_data_out(46), S0=>nx36231);
   ix15784 : mux21_ni port map ( Y=>nx15783, A0=>label_3_output(13), A1=>
      label_3_input_13, S0=>nx36269);
   ix3493 : mux21_ni port map ( Y=>nx3492, A0=>nx3488, A1=>
      label_3_input_state_machine_13, S0=>nx35949);
   ix15774 : mux21_ni port map ( Y=>nx15773, A0=>
      label_3_input_state_machine_13, A1=>mdr_data_out(45), S0=>nx36231);
   ix15744 : mux21_ni port map ( Y=>nx15743, A0=>label_3_output(11), A1=>
      label_3_input_11, S0=>nx36269);
   ix3429 : mux21_ni port map ( Y=>nx3428, A0=>nx3424, A1=>
      label_3_input_state_machine_11, S0=>nx35949);
   ix15734 : mux21_ni port map ( Y=>nx15733, A0=>
      label_3_input_state_machine_11, A1=>mdr_data_out(43), S0=>nx36231);
   ix15704 : mux21_ni port map ( Y=>nx15703, A0=>label_3_output(9), A1=>
      label_3_input_9, S0=>nx36269);
   ix3365 : mux21_ni port map ( Y=>nx3364, A0=>nx3360, A1=>
      label_3_input_state_machine_9, S0=>nx35947);
   ix15694 : mux21_ni port map ( Y=>nx15693, A0=>
      label_3_input_state_machine_9, A1=>mdr_data_out(41), S0=>nx36231);
   ix15664 : mux21_ni port map ( Y=>nx15663, A0=>label_3_output(7), A1=>
      label_3_input_7, S0=>nx36269);
   ix3301 : mux21_ni port map ( Y=>nx3300, A0=>nx3296, A1=>
      label_3_input_state_machine_7, S0=>nx35947);
   ix15654 : mux21_ni port map ( Y=>nx15653, A0=>
      label_3_input_state_machine_7, A1=>mdr_data_out(39), S0=>nx36233);
   ix15624 : mux21_ni port map ( Y=>nx15623, A0=>label_3_output(5), A1=>
      label_3_input_5, S0=>nx36271);
   ix3237 : mux21_ni port map ( Y=>nx3236, A0=>nx3232, A1=>
      label_3_input_state_machine_5, S0=>nx35169);
   ix15614 : mux21_ni port map ( Y=>nx15613, A0=>
      label_3_input_state_machine_5, A1=>mdr_data_out(37), S0=>nx36233);
   ix15584 : mux21_ni port map ( Y=>nx15583, A0=>label_3_output(3), A1=>
      label_3_input_3, S0=>nx36271);
   ix3173 : mux21_ni port map ( Y=>nx3172, A0=>nx3168, A1=>
      label_3_input_state_machine_3, S0=>nx35169);
   ix15574 : mux21_ni port map ( Y=>nx15573, A0=>
      label_3_input_state_machine_3, A1=>mdr_data_out(35), S0=>nx36233);
   ix15544 : mux21_ni port map ( Y=>nx15543, A0=>label_3_output(1), A1=>
      label_3_input_1, S0=>nx36271);
   ix3109 : mux21_ni port map ( Y=>nx3108, A0=>nx3104, A1=>
      label_3_input_state_machine_1, S0=>nx35169);
   ix15534 : mux21_ni port map ( Y=>nx15533, A0=>
      label_3_input_state_machine_1, A1=>mdr_data_out(33), S0=>nx36233);
   ix32765 : xnor2 port map ( Y=>nx32764, A0=>nx29051, A1=>nx32774);
   ix15564 : mux21_ni port map ( Y=>nx15563, A0=>label_3_output(2), A1=>
      label_3_input_2, S0=>nx36271);
   ix3141 : mux21_ni port map ( Y=>nx3140, A0=>nx3136, A1=>
      label_3_input_state_machine_2, S0=>nx35169);
   ix15554 : mux21_ni port map ( Y=>nx15553, A0=>
      label_3_input_state_machine_2, A1=>mdr_data_out(34), S0=>nx36233);
   ix32780 : xnor2 port map ( Y=>nx32779, A0=>nx29049, A1=>nx32789);
   ix15604 : mux21_ni port map ( Y=>nx15603, A0=>label_3_output(4), A1=>
      label_3_input_4, S0=>nx36271);
   ix3205 : mux21_ni port map ( Y=>nx3204, A0=>nx3200, A1=>
      label_3_input_state_machine_4, S0=>nx35169);
   ix15594 : mux21_ni port map ( Y=>nx15593, A0=>
      label_3_input_state_machine_4, A1=>mdr_data_out(36), S0=>nx36233);
   ix32795 : xnor2 port map ( Y=>nx32794, A0=>nx29047, A1=>nx32804);
   ix15644 : mux21_ni port map ( Y=>nx15643, A0=>label_3_output(6), A1=>
      label_3_input_6, S0=>nx36271);
   ix3269 : mux21_ni port map ( Y=>nx3268, A0=>nx3264, A1=>
      label_3_input_state_machine_6, S0=>nx35169);
   ix15634 : mux21_ni port map ( Y=>nx15633, A0=>
      label_3_input_state_machine_6, A1=>mdr_data_out(38), S0=>nx36233);
   ix32810 : xnor2 port map ( Y=>nx32809, A0=>nx29045, A1=>nx32819);
   ix15684 : mux21_ni port map ( Y=>nx15683, A0=>label_3_output(8), A1=>
      label_3_input_8, S0=>nx36271);
   ix3333 : mux21_ni port map ( Y=>nx3332, A0=>nx3328, A1=>
      label_3_input_state_machine_8, S0=>nx35169);
   ix15674 : mux21_ni port map ( Y=>nx15673, A0=>
      label_3_input_state_machine_8, A1=>mdr_data_out(40), S0=>nx36235);
   ix32825 : xnor2 port map ( Y=>nx32824, A0=>nx29043, A1=>nx32834);
   ix15724 : mux21_ni port map ( Y=>nx15723, A0=>label_3_output(10), A1=>
      label_3_input_10, S0=>nx36273);
   ix3397 : mux21_ni port map ( Y=>nx3396, A0=>nx3392, A1=>
      label_3_input_state_machine_10, S0=>nx35949);
   ix15714 : mux21_ni port map ( Y=>nx15713, A0=>
      label_3_input_state_machine_10, A1=>mdr_data_out(42), S0=>nx36235);
   ix32840 : xnor2 port map ( Y=>nx32839, A0=>nx29041, A1=>nx32849);
   ix15764 : mux21_ni port map ( Y=>nx15763, A0=>label_3_output(12), A1=>
      label_3_input_12, S0=>nx36273);
   ix3461 : mux21_ni port map ( Y=>nx3460, A0=>nx3456, A1=>
      label_3_input_state_machine_12, S0=>nx35949);
   ix15754 : mux21_ni port map ( Y=>nx15753, A0=>
      label_3_input_state_machine_12, A1=>mdr_data_out(44), S0=>nx36235);
   ix32855 : xnor2 port map ( Y=>nx32854, A0=>nx29039, A1=>nx32856);
   ix21664 : ao32 port map ( Y=>nx21663, A0=>nx35961, A1=>nx35653, A2=>
      nx36293, B0=>max_calc_ans3_14, B1=>nx35877);
   ix32860 : mux21 port map ( Y=>nx35653, A0=>nx29942, A1=>nx30132, S0=>
      nx35887);
   ix15909 : xnor2 port map ( Y=>nx15908, A0=>nx32472, A1=>nx32669);
   ix32866 : xnor2 port map ( Y=>nx32865, A0=>nx32869, A1=>
      max_calc_comparator_second_inp1_13);
   ix15935 : mux21_ni port map ( Y=>nx15934, A0=>max_calc_ans4_13, A1=>
      label_4_output(13), S0=>nx35979);
   ix23724 : ao32 port map ( Y=>nx23723, A0=>nx35961, A1=>nx35655, A2=>
      nx36293, B0=>max_calc_ans4_13, B1=>nx35877);
   ix32877 : mux21 port map ( Y=>nx35655, A0=>nx32252, A1=>nx32256, S0=>
      nx35893);
   ix15971 : mux21_ni port map ( Y=>nx15970, A0=>max_calc_ans3_13, A1=>
      label_3_output(13), S0=>nx35979);
   ix23744 : ao32 port map ( Y=>nx23743, A0=>nx35961, A1=>nx35657, A2=>
      nx36293, B0=>max_calc_ans3_13, B1=>nx35877);
   ix32889 : mux21 port map ( Y=>nx35657, A0=>nx30325, A1=>nx30329, S0=>
      nx35887);
   ix16009 : mux21 port map ( Y=>nx16008, A0=>nx32904, A1=>nx32653, S0=>
      nx35979);
   ix23764 : ao32 port map ( Y=>nx23763, A0=>nx35961, A1=>nx35659, A2=>
      nx36293, B0=>max_calc_ans4_12, B1=>nx35877);
   ix32903 : mux21 port map ( Y=>nx35659, A0=>nx32263, A1=>nx32270, S0=>
      nx35893);
   ix16045 : mux21 port map ( Y=>nx16044, A0=>nx32917, A1=>nx32849, S0=>
      nx35981);
   ix23784 : ao32 port map ( Y=>nx23783, A0=>nx35961, A1=>nx35661, A2=>
      nx36293, B0=>max_calc_ans3_12, B1=>nx35879);
   ix32916 : mux21 port map ( Y=>nx35661, A0=>nx30336, A1=>nx30343, S0=>
      nx35887);
   ix16057 : xnor2 port map ( Y=>nx16056, A0=>nx32894, A1=>nx32908);
   ix32922 : xnor2 port map ( Y=>nx32921, A0=>nx32925, A1=>
      max_calc_comparator_second_inp1_11);
   ix16083 : mux21_ni port map ( Y=>nx16082, A0=>max_calc_ans4_11, A1=>
      label_4_output(11), S0=>nx35981);
   ix23804 : ao32 port map ( Y=>nx23803, A0=>nx35963, A1=>nx35663, A2=>
      nx36293, B0=>max_calc_ans4_11, B1=>nx35879);
   ix32933 : mux21 port map ( Y=>nx35663, A0=>nx32280, A1=>nx32284, S0=>
      nx35893);
   ix16119 : mux21_ni port map ( Y=>nx16118, A0=>max_calc_ans3_11, A1=>
      label_3_output(11), S0=>nx35981);
   ix23824 : ao32 port map ( Y=>nx23823, A0=>nx35963, A1=>nx35665, A2=>
      nx36293, B0=>max_calc_ans3_11, B1=>nx35879);
   ix32945 : mux21 port map ( Y=>nx35665, A0=>nx30353, A1=>nx30357, S0=>
      nx35887);
   ix16157 : mux21 port map ( Y=>nx16156, A0=>nx32960, A1=>nx32638, S0=>
      nx35981);
   ix23844 : ao32 port map ( Y=>nx23843, A0=>nx35963, A1=>nx35667, A2=>
      nx36295, B0=>max_calc_ans4_10, B1=>nx35879);
   ix32959 : mux21 port map ( Y=>nx35667, A0=>nx32291, A1=>nx32298, S0=>
      nx35893);
   ix16193 : mux21 port map ( Y=>nx16192, A0=>nx32973, A1=>nx32834, S0=>
      nx35981);
   ix23864 : ao32 port map ( Y=>nx23863, A0=>nx35963, A1=>nx35669, A2=>
      nx36295, B0=>max_calc_ans3_10, B1=>nx35879);
   ix32972 : mux21 port map ( Y=>nx35669, A0=>nx30364, A1=>nx30371, S0=>
      nx35887);
   ix16205 : xnor2 port map ( Y=>nx16204, A0=>nx32950, A1=>nx32964);
   ix32978 : xnor2 port map ( Y=>nx32977, A0=>nx32981, A1=>
      max_calc_comparator_second_inp1_9);
   ix16231 : mux21_ni port map ( Y=>nx16230, A0=>max_calc_ans4_9, A1=>
      label_4_output(9), S0=>nx35981);
   ix23884 : ao32 port map ( Y=>nx23883, A0=>nx35963, A1=>nx35671, A2=>
      nx36295, B0=>max_calc_ans4_9, B1=>nx35879);
   ix32989 : mux21 port map ( Y=>nx35671, A0=>nx32308, A1=>nx32312, S0=>
      nx35893);
   ix16267 : mux21_ni port map ( Y=>nx16266, A0=>max_calc_ans3_9, A1=>
      label_3_output(9), S0=>nx35981);
   ix23904 : ao32 port map ( Y=>nx23903, A0=>nx35963, A1=>nx35673, A2=>
      nx36295, B0=>max_calc_ans3_9, B1=>nx35879);
   ix33001 : mux21 port map ( Y=>nx35673, A0=>nx30381, A1=>nx30385, S0=>
      nx35887);
   ix16305 : mux21 port map ( Y=>nx16304, A0=>nx33016, A1=>nx32623, S0=>
      nx35983);
   ix23924 : ao32 port map ( Y=>nx23923, A0=>nx35963, A1=>nx35675, A2=>
      nx36295, B0=>max_calc_ans4_8, B1=>nx35881);
   ix33015 : mux21 port map ( Y=>nx35675, A0=>nx32319, A1=>nx32326, S0=>
      nx35895);
   ix16341 : mux21 port map ( Y=>nx16340, A0=>nx33029, A1=>nx32819, S0=>
      nx35983);
   ix23944 : ao32 port map ( Y=>nx23943, A0=>nx35183, A1=>nx35677, A2=>
      nx36295, B0=>max_calc_ans3_8, B1=>nx35881);
   ix33028 : mux21 port map ( Y=>nx35677, A0=>nx30392, A1=>nx30399, S0=>
      nx35889);
   ix16353 : xnor2 port map ( Y=>nx16352, A0=>nx33006, A1=>nx33020);
   ix33034 : xnor2 port map ( Y=>nx33033, A0=>nx33037, A1=>
      max_calc_comparator_second_inp1_7);
   ix16379 : mux21_ni port map ( Y=>nx16378, A0=>max_calc_ans4_7, A1=>
      label_4_output(7), S0=>nx35983);
   ix23964 : ao32 port map ( Y=>nx23963, A0=>nx35183, A1=>nx35679, A2=>
      nx36295, B0=>max_calc_ans4_7, B1=>nx35881);
   ix33045 : mux21 port map ( Y=>nx35679, A0=>nx32336, A1=>nx32340, S0=>
      nx35895);
   ix16415 : mux21_ni port map ( Y=>nx16414, A0=>max_calc_ans3_7, A1=>
      label_3_output(7), S0=>nx35983);
   ix23984 : ao32 port map ( Y=>nx23983, A0=>nx35183, A1=>nx35681, A2=>
      nx36297, B0=>max_calc_ans3_7, B1=>nx35881);
   ix33057 : mux21 port map ( Y=>nx35681, A0=>nx30409, A1=>nx30413, S0=>
      nx35889);
   ix16453 : mux21 port map ( Y=>nx16452, A0=>nx33072, A1=>nx32608, S0=>
      nx35983);
   ix24004 : ao32 port map ( Y=>nx24003, A0=>nx35965, A1=>nx35683, A2=>
      nx36297, B0=>max_calc_ans4_6, B1=>nx35881);
   ix33071 : mux21 port map ( Y=>nx35683, A0=>nx32347, A1=>nx32354, S0=>
      nx35895);
   ix16489 : mux21 port map ( Y=>nx16488, A0=>nx33085, A1=>nx32804, S0=>
      nx35983);
   ix24024 : ao32 port map ( Y=>nx24023, A0=>nx35965, A1=>nx35685, A2=>
      nx36297, B0=>max_calc_ans3_6, B1=>nx35881);
   ix33084 : mux21 port map ( Y=>nx35685, A0=>nx30420, A1=>nx30427, S0=>
      nx35889);
   ix16501 : xnor2 port map ( Y=>nx16500, A0=>nx33062, A1=>nx33076);
   ix33090 : xnor2 port map ( Y=>nx33089, A0=>nx33093, A1=>
      max_calc_comparator_second_inp1_5);
   ix16527 : mux21_ni port map ( Y=>nx16526, A0=>max_calc_ans4_5, A1=>
      label_4_output(5), S0=>nx35983);
   ix24044 : ao32 port map ( Y=>nx24043, A0=>nx35965, A1=>nx35687, A2=>
      nx36297, B0=>max_calc_ans4_5, B1=>nx35881);
   ix33101 : mux21 port map ( Y=>nx35687, A0=>nx32364, A1=>nx32368, S0=>
      nx35895);
   ix16563 : mux21_ni port map ( Y=>nx16562, A0=>max_calc_ans3_5, A1=>
      label_3_output(5), S0=>nx35985);
   ix24064 : ao32 port map ( Y=>nx24063, A0=>nx35965, A1=>nx35689, A2=>
      nx36297, B0=>max_calc_ans3_5, B1=>nx35883);
   ix33113 : mux21 port map ( Y=>nx35689, A0=>nx30437, A1=>nx30441, S0=>
      nx35889);
   ix16601 : mux21 port map ( Y=>nx16600, A0=>nx33128, A1=>nx32593, S0=>
      nx35985);
   ix24084 : ao32 port map ( Y=>nx24083, A0=>nx35965, A1=>nx35691, A2=>
      nx36297, B0=>max_calc_ans4_4, B1=>nx35883);
   ix33127 : mux21 port map ( Y=>nx35691, A0=>nx32375, A1=>nx32382, S0=>
      nx35895);
   ix16637 : mux21 port map ( Y=>nx16636, A0=>nx33141, A1=>nx32789, S0=>
      nx35985);
   ix24104 : ao32 port map ( Y=>nx24103, A0=>nx35965, A1=>nx35693, A2=>
      nx36297, B0=>max_calc_ans3_4, B1=>nx35883);
   ix33140 : mux21 port map ( Y=>nx35693, A0=>nx30448, A1=>nx30455, S0=>
      nx35889);
   ix16649 : xnor2 port map ( Y=>nx16648, A0=>nx33118, A1=>nx33132);
   ix33146 : xnor2 port map ( Y=>nx33145, A0=>nx33149, A1=>
      max_calc_comparator_second_inp1_3);
   ix16675 : mux21_ni port map ( Y=>nx16674, A0=>max_calc_ans4_3, A1=>
      label_4_output(3), S0=>nx35985);
   ix24124 : ao32 port map ( Y=>nx24123, A0=>nx35967, A1=>nx35695, A2=>
      nx36393, B0=>max_calc_ans4_3, B1=>nx35883);
   ix33157 : mux21 port map ( Y=>nx35695, A0=>nx32392, A1=>nx32396, S0=>
      nx35895);
   ix16711 : mux21_ni port map ( Y=>nx16710, A0=>max_calc_ans3_3, A1=>
      label_3_output(3), S0=>nx35985);
   ix24144 : ao32 port map ( Y=>nx24143, A0=>nx35967, A1=>nx35697, A2=>
      nx36393, B0=>max_calc_ans3_3, B1=>nx35883);
   ix33169 : mux21 port map ( Y=>nx35697, A0=>nx30465, A1=>nx30469, S0=>
      nx35889);
   ix16749 : mux21 port map ( Y=>nx16748, A0=>nx33184, A1=>nx32578, S0=>
      nx35985);
   ix24164 : ao32 port map ( Y=>nx24163, A0=>nx35967, A1=>nx35699, A2=>
      nx36393, B0=>max_calc_ans4_2, B1=>nx35883);
   ix33183 : mux21 port map ( Y=>nx35699, A0=>nx32403, A1=>nx32410, S0=>
      nx35895);
   ix16785 : mux21 port map ( Y=>nx16784, A0=>nx33197, A1=>nx32774, S0=>
      nx35985);
   ix24184 : ao32 port map ( Y=>nx24183, A0=>nx35967, A1=>nx35701, A2=>
      nx36393, B0=>max_calc_ans3_2, B1=>nx35883);
   ix33196 : mux21 port map ( Y=>nx35701, A0=>nx30476, A1=>nx30483, S0=>
      nx35889);
   ix16797 : xnor2 port map ( Y=>nx16796, A0=>nx33174, A1=>nx33188);
   ix16823 : mux21_ni port map ( Y=>nx16822, A0=>max_calc_ans4_1, A1=>
      label_4_output(1), S0=>nx35187);
   ix24204 : ao32 port map ( Y=>nx24203, A0=>nx35967, A1=>nx35703, A2=>
      nx36393, B0=>max_calc_ans4_1, B1=>nx35885);
   ix33211 : mux21 port map ( Y=>nx35703, A0=>nx32418, A1=>nx32422, S0=>
      nx35897);
   ix16859 : mux21_ni port map ( Y=>nx16858, A0=>max_calc_ans3_1, A1=>
      label_3_output(1), S0=>nx35987);
   ix24224 : ao32 port map ( Y=>nx24223, A0=>nx35967, A1=>nx35705, A2=>
      nx36393, B0=>max_calc_ans3_1, B1=>nx35885);
   ix33223 : mux21 port map ( Y=>nx35705, A0=>nx30491, A1=>nx30495, S0=>
      nx35891);
   ix16871 : xnor2 port map ( Y=>nx16870, A0=>nx33203, A1=>nx33214);
   ix17137 : xnor2 port map ( Y=>nx17136, A0=>nx33232, A1=>nx33257);
   ix17089 : mux21_ni port map ( Y=>nx17088, A0=>max_calc_ans4_15, A1=>
      label_4_output(15), S0=>nx35987);
   ix14964 : mux21_ni port map ( Y=>nx14963, A0=>label_4_output(15), A1=>
      label_4_input_15, S0=>nx36273);
   ix2213 : mux21_ni port map ( Y=>nx2212, A0=>nx2208, A1=>
      label_4_input_state_machine_15, S0=>nx35949);
   ix14124 : mux21_ni port map ( Y=>nx14123, A0=>
      label_4_input_state_machine_15, A1=>mdr_data_out(63), S0=>nx36235);
   ix33247 : xor2 port map ( Y=>nx33246, A0=>nx30966, A1=>label_4_output(15)
   );
   ix24284 : ao32 port map ( Y=>nx24283, A0=>nx35967, A1=>nx35707, A2=>
      nx36393, B0=>max_calc_ans4_15, B1=>nx35885);
   ix33252 : mux21 port map ( Y=>nx35707, A0=>nx32433, A1=>nx32451, S0=>
      nx35897);
   ix17125 : mux21_ni port map ( Y=>nx17124, A0=>max_calc_ans3_15, A1=>
      label_3_output(15), S0=>nx35987);
   ix15814 : mux21_ni port map ( Y=>nx15813, A0=>label_3_output(15), A1=>
      label_3_input_15, S0=>nx36273);
   ix3551 : mux21_ni port map ( Y=>nx3550, A0=>nx3546, A1=>
      label_3_input_state_machine_15, S0=>nx35949);
   ix14974 : mux21_ni port map ( Y=>nx14973, A0=>
      label_3_input_state_machine_15, A1=>mdr_data_out(47), S0=>nx36235);
   ix33272 : xor2 port map ( Y=>nx33271, A0=>nx29037, A1=>label_3_output(15)
   );
   ix24304 : ao32 port map ( Y=>nx24303, A0=>nx35969, A1=>nx35709, A2=>
      nx35749, B0=>max_calc_ans3_15, B1=>nx35885);
   ix33277 : mux21 port map ( Y=>nx35709, A0=>nx30506, A1=>nx30524, S0=>
      nx35891);
   ix18889 : mux21_ni port map ( Y=>nx18888, A0=>max_calc_ans8_0, A1=>
      max_calc_ans7_0, S0=>nx35987);
   ix25464 : mux21_ni port map ( Y=>nx25463, A0=>max_calc_ans7_0, A1=>
      nx18854, S0=>nx36021);
   ix25454 : mux21_ni port map ( Y=>nx25453, A0=>nx13121, A1=>
      max_calc_ans8_0, S0=>nx35869);
   ix24394 : mux21_ni port map ( Y=>nx24393, A0=>
      max_calc_comparator_first_inp2_14, A1=>nx17248, S0=>nx36281);
   ix17249 : mux21_ni port map ( Y=>nx17248, A0=>nx17244, A1=>nx17156, S0=>
      nx35969);
   ix17157 : mux21_ni port map ( Y=>nx17156, A0=>max_calc_ans2_14, A1=>
      label_2_output(14), S0=>nx35987);
   ix16654 : mux21_ni port map ( Y=>nx16653, A0=>label_2_output(14), A1=>
      label_2_input_14, S0=>nx36273);
   ix4863 : mux21_ni port map ( Y=>nx4862, A0=>nx4858, A1=>
      label_2_input_state_machine_14, S0=>nx35951);
   ix16644 : mux21_ni port map ( Y=>nx16643, A0=>
      label_2_input_state_machine_14, A1=>mdr_data_out(30), S0=>nx36235);
   ix16634 : mux21_ni port map ( Y=>nx16633, A0=>label_2_output(13), A1=>
      label_2_input_13, S0=>nx36273);
   ix4831 : mux21_ni port map ( Y=>nx4830, A0=>nx4826, A1=>
      label_2_input_state_machine_13, S0=>nx35951);
   ix16624 : mux21_ni port map ( Y=>nx16623, A0=>
      label_2_input_state_machine_13, A1=>mdr_data_out(29), S0=>nx36235);
   ix16594 : mux21_ni port map ( Y=>nx16593, A0=>label_2_output(11), A1=>
      label_2_input_11, S0=>nx36273);
   ix4767 : mux21_ni port map ( Y=>nx4766, A0=>nx4762, A1=>
      label_2_input_state_machine_11, S0=>nx35951);
   ix16584 : mux21_ni port map ( Y=>nx16583, A0=>
      label_2_input_state_machine_11, A1=>mdr_data_out(27), S0=>nx35599);
   ix16554 : mux21_ni port map ( Y=>nx16553, A0=>label_2_output(9), A1=>
      label_2_input_9, S0=>nx36275);
   ix4703 : mux21_ni port map ( Y=>nx4702, A0=>nx4698, A1=>
      label_2_input_state_machine_9, S0=>nx35951);
   ix16544 : mux21_ni port map ( Y=>nx16543, A0=>
      label_2_input_state_machine_9, A1=>mdr_data_out(25), S0=>nx35599);
   ix16514 : mux21_ni port map ( Y=>nx16513, A0=>label_2_output(7), A1=>
      label_2_input_7, S0=>nx36275);
   ix4639 : mux21_ni port map ( Y=>nx4638, A0=>nx4634, A1=>
      label_2_input_state_machine_7, S0=>nx35951);
   ix16504 : mux21_ni port map ( Y=>nx16503, A0=>
      label_2_input_state_machine_7, A1=>mdr_data_out(23), S0=>nx35599);
   ix16474 : mux21_ni port map ( Y=>nx16473, A0=>label_2_output(5), A1=>
      label_2_input_5, S0=>nx36275);
   ix4575 : mux21_ni port map ( Y=>nx4574, A0=>nx4570, A1=>
      label_2_input_state_machine_5, S0=>nx35951);
   ix16464 : mux21_ni port map ( Y=>nx16463, A0=>
      label_2_input_state_machine_5, A1=>mdr_data_out(21), S0=>nx35599);
   ix16434 : mux21_ni port map ( Y=>nx16433, A0=>label_2_output(3), A1=>
      label_2_input_3, S0=>nx36275);
   ix4511 : mux21_ni port map ( Y=>nx4510, A0=>nx4506, A1=>
      label_2_input_state_machine_3, S0=>nx35951);
   ix16424 : mux21_ni port map ( Y=>nx16423, A0=>
      label_2_input_state_machine_3, A1=>mdr_data_out(19), S0=>nx35599);
   ix16394 : mux21_ni port map ( Y=>nx16393, A0=>label_2_output(1), A1=>
      label_2_input_1, S0=>nx36275);
   ix4447 : mux21_ni port map ( Y=>nx4446, A0=>nx4442, A1=>
      label_2_input_state_machine_1, S0=>nx35953);
   ix16384 : mux21_ni port map ( Y=>nx16383, A0=>
      label_2_input_state_machine_1, A1=>mdr_data_out(17), S0=>nx35599);
   ix33388 : xnor2 port map ( Y=>nx33387, A0=>nx28608, A1=>nx33397);
   ix16414 : mux21_ni port map ( Y=>nx16413, A0=>label_2_output(2), A1=>
      label_2_input_2, S0=>nx36275);
   ix4479 : mux21_ni port map ( Y=>nx4478, A0=>nx4474, A1=>
      label_2_input_state_machine_2, S0=>nx35953);
   ix16404 : mux21_ni port map ( Y=>nx16403, A0=>
      label_2_input_state_machine_2, A1=>mdr_data_out(18), S0=>nx35599);
   ix33403 : xnor2 port map ( Y=>nx33402, A0=>nx28606, A1=>nx33412);
   ix16454 : mux21_ni port map ( Y=>nx16453, A0=>label_2_output(4), A1=>
      label_2_input_4, S0=>nx36275);
   ix4543 : mux21_ni port map ( Y=>nx4542, A0=>nx4538, A1=>
      label_2_input_state_machine_4, S0=>nx35953);
   ix16444 : mux21_ni port map ( Y=>nx16443, A0=>
      label_2_input_state_machine_4, A1=>mdr_data_out(20), S0=>nx36237);
   ix33418 : xnor2 port map ( Y=>nx33417, A0=>nx28604, A1=>nx33427);
   ix16494 : mux21_ni port map ( Y=>nx16493, A0=>label_2_output(6), A1=>
      label_2_input_6, S0=>nx35607);
   ix4607 : mux21_ni port map ( Y=>nx4606, A0=>nx4602, A1=>
      label_2_input_state_machine_6, S0=>nx35953);
   ix16484 : mux21_ni port map ( Y=>nx16483, A0=>
      label_2_input_state_machine_6, A1=>mdr_data_out(22), S0=>nx36237);
   ix33433 : xnor2 port map ( Y=>nx33432, A0=>nx28602, A1=>nx33442);
   ix16534 : mux21_ni port map ( Y=>nx16533, A0=>label_2_output(8), A1=>
      label_2_input_8, S0=>nx35607);
   ix4671 : mux21_ni port map ( Y=>nx4670, A0=>nx4666, A1=>
      label_2_input_state_machine_8, S0=>nx35953);
   ix16524 : mux21_ni port map ( Y=>nx16523, A0=>
      label_2_input_state_machine_8, A1=>mdr_data_out(24), S0=>nx36237);
   ix33448 : xnor2 port map ( Y=>nx33447, A0=>nx28600, A1=>nx33457);
   ix16574 : mux21_ni port map ( Y=>nx16573, A0=>label_2_output(10), A1=>
      label_2_input_10, S0=>nx35607);
   ix4735 : mux21_ni port map ( Y=>nx4734, A0=>nx4730, A1=>
      label_2_input_state_machine_10, S0=>nx35953);
   ix16564 : mux21_ni port map ( Y=>nx16563, A0=>
      label_2_input_state_machine_10, A1=>mdr_data_out(26), S0=>nx36237);
   ix33463 : xnor2 port map ( Y=>nx33462, A0=>nx28598, A1=>nx33472);
   ix16614 : mux21_ni port map ( Y=>nx16613, A0=>label_2_output(12), A1=>
      label_2_input_12, S0=>nx35607);
   ix4799 : mux21_ni port map ( Y=>nx4798, A0=>nx4794, A1=>
      label_2_input_state_machine_12, S0=>nx35953);
   ix16604 : mux21_ni port map ( Y=>nx16603, A0=>
      label_2_input_state_machine_12, A1=>mdr_data_out(28), S0=>nx36237);
   ix33478 : xnor2 port map ( Y=>nx33477, A0=>nx28596, A1=>nx33479);
   ix24324 : mux21_ni port map ( Y=>nx24323, A0=>nx17146, A1=>
      max_calc_ans2_14, S0=>nx35851);
   ix17147 : mux21 port map ( Y=>nx17146, A0=>nx32472, A1=>nx32669, S0=>
      nx35899);
   ix17245 : mux21_ni port map ( Y=>nx17244, A0=>max_calc_ans8_14, A1=>
      max_calc_ans7_14, S0=>nx35987);
   ix24384 : mux21_ni port map ( Y=>nx24383, A0=>max_calc_ans7_14, A1=>
      nx17146, S0=>nx36021);
   ix24374 : mux21_ni port map ( Y=>nx24373, A0=>nx13371, A1=>
      max_calc_ans8_14, S0=>nx35869);
   ix17225 : mux21_ni port map ( Y=>nx13371, A0=>
      max_calc_comparator_first_inp2_14, A1=>
      max_calc_comparator_first_inp1_14, S0=>nx35905);
   ix24364 : mux21_ni port map ( Y=>nx24363, A0=>
      max_calc_comparator_first_inp1_14, A1=>nx17210, S0=>nx36281);
   ix17211 : mux21_ni port map ( Y=>nx17210, A0=>nx17206, A1=>nx17174, S0=>
      nx35969);
   ix17175 : mux21_ni port map ( Y=>nx17174, A0=>max_calc_ans1_14, A1=>
      label_1_output(14), S0=>nx35989);
   ix17504 : mux21_ni port map ( Y=>nx17503, A0=>label_1_output(14), A1=>
      label_1_input_14, S0=>nx36277);
   ix6201 : mux21_ni port map ( Y=>nx6200, A0=>nx6196, A1=>
      label_1_input_state_machine_14, S0=>nx35955);
   ix17494 : mux21_ni port map ( Y=>nx17493, A0=>
      label_1_input_state_machine_14, A1=>mdr_data_out(14), S0=>nx36237);
   ix17484 : mux21_ni port map ( Y=>nx17483, A0=>label_1_output(13), A1=>
      label_1_input_13, S0=>nx36277);
   ix6169 : mux21_ni port map ( Y=>nx6168, A0=>nx6164, A1=>
      label_1_input_state_machine_13, S0=>nx35955);
   ix17474 : mux21_ni port map ( Y=>nx17473, A0=>
      label_1_input_state_machine_13, A1=>mdr_data_out(13), S0=>nx36237);
   ix17444 : mux21_ni port map ( Y=>nx17443, A0=>label_1_output(11), A1=>
      label_1_input_11, S0=>nx36279);
   ix6105 : mux21_ni port map ( Y=>nx6104, A0=>nx6100, A1=>
      label_1_input_state_machine_11, S0=>nx35955);
   ix17434 : mux21_ni port map ( Y=>nx17433, A0=>
      label_1_input_state_machine_11, A1=>mdr_data_out(11), S0=>nx36239);
   ix17404 : mux21_ni port map ( Y=>nx17403, A0=>label_1_output(9), A1=>
      label_1_input_9, S0=>nx36279);
   ix6041 : mux21_ni port map ( Y=>nx6040, A0=>nx6036, A1=>
      label_1_input_state_machine_9, S0=>nx35955);
   ix17394 : mux21_ni port map ( Y=>nx17393, A0=>
      label_1_input_state_machine_9, A1=>mdr_data_out(9), S0=>nx36239);
   ix17364 : mux21_ni port map ( Y=>nx17363, A0=>label_1_output(7), A1=>
      label_1_input_7, S0=>nx36279);
   ix5977 : mux21_ni port map ( Y=>nx5976, A0=>nx5972, A1=>
      label_1_input_state_machine_7, S0=>nx35955);
   ix17354 : mux21_ni port map ( Y=>nx17353, A0=>
      label_1_input_state_machine_7, A1=>mdr_data_out(7), S0=>nx36239);
   ix17324 : mux21_ni port map ( Y=>nx17323, A0=>label_1_output(5), A1=>
      label_1_input_5, S0=>nx36279);
   ix5913 : mux21_ni port map ( Y=>nx5912, A0=>nx5908, A1=>
      label_1_input_state_machine_5, S0=>nx35955);
   ix17314 : mux21_ni port map ( Y=>nx17313, A0=>
      label_1_input_state_machine_5, A1=>mdr_data_out(5), S0=>nx36239);
   ix17284 : mux21_ni port map ( Y=>nx17283, A0=>label_1_output(3), A1=>
      label_1_input_3, S0=>nx35607);
   ix5849 : mux21_ni port map ( Y=>nx5848, A0=>nx5844, A1=>
      label_1_input_state_machine_3, S0=>nx35955);
   ix17274 : mux21_ni port map ( Y=>nx17273, A0=>
      label_1_input_state_machine_3, A1=>mdr_data_out(3), S0=>nx36239);
   ix17244 : mux21_ni port map ( Y=>nx17243, A0=>label_1_output(1), A1=>
      label_1_input_1, S0=>nx35607);
   ix5785 : mux21_ni port map ( Y=>nx5784, A0=>nx5780, A1=>
      label_1_input_state_machine_1, S0=>nx35957);
   ix17234 : mux21_ni port map ( Y=>nx17233, A0=>
      label_1_input_state_machine_1, A1=>mdr_data_out(1), S0=>nx36239);
   ix33586 : xnor2 port map ( Y=>nx33585, A0=>nx26648, A1=>nx33595);
   ix17264 : mux21_ni port map ( Y=>nx17263, A0=>label_1_output(2), A1=>
      label_1_input_2, S0=>nx35607);
   ix5817 : mux21_ni port map ( Y=>nx5816, A0=>nx5812, A1=>
      label_1_input_state_machine_2, S0=>nx35957);
   ix17254 : mux21_ni port map ( Y=>nx17253, A0=>
      label_1_input_state_machine_2, A1=>mdr_data_out(2), S0=>nx36239);
   ix33601 : xnor2 port map ( Y=>nx33600, A0=>nx26646, A1=>nx33610);
   ix17304 : mux21_ni port map ( Y=>nx17303, A0=>label_1_output(4), A1=>
      label_1_input_4, S0=>nx36279);
   ix5881 : mux21_ni port map ( Y=>nx5880, A0=>nx5876, A1=>
      label_1_input_state_machine_4, S0=>nx35957);
   ix17294 : mux21_ni port map ( Y=>nx17293, A0=>
      label_1_input_state_machine_4, A1=>mdr_data_out(4), S0=>nx35601);
   ix33616 : xnor2 port map ( Y=>nx33615, A0=>nx26644, A1=>nx33625);
   ix17344 : mux21_ni port map ( Y=>nx17343, A0=>label_1_output(6), A1=>
      label_1_input_6, S0=>nx36279);
   ix5945 : mux21_ni port map ( Y=>nx5944, A0=>nx5940, A1=>
      label_1_input_state_machine_6, S0=>nx35957);
   ix17334 : mux21_ni port map ( Y=>nx17333, A0=>
      label_1_input_state_machine_6, A1=>mdr_data_out(6), S0=>nx35601);
   ix33631 : xnor2 port map ( Y=>nx33630, A0=>nx26642, A1=>nx33640);
   ix17384 : mux21_ni port map ( Y=>nx17383, A0=>label_1_output(8), A1=>
      label_1_input_8, S0=>nx36279);
   ix6009 : mux21_ni port map ( Y=>nx6008, A0=>nx6004, A1=>
      label_1_input_state_machine_8, S0=>nx35957);
   ix17374 : mux21_ni port map ( Y=>nx17373, A0=>
      label_1_input_state_machine_8, A1=>mdr_data_out(8), S0=>nx35601);
   ix33646 : xnor2 port map ( Y=>nx33645, A0=>nx26640, A1=>nx33655);
   ix17424 : mux21_ni port map ( Y=>nx17423, A0=>label_1_output(10), A1=>
      label_1_input_10, S0=>nx35609);
   ix6073 : mux21_ni port map ( Y=>nx6072, A0=>nx6068, A1=>
      label_1_input_state_machine_10, S0=>nx35957);
   ix17414 : mux21_ni port map ( Y=>nx17413, A0=>
      label_1_input_state_machine_10, A1=>mdr_data_out(10), S0=>nx35601);
   ix33661 : xnor2 port map ( Y=>nx33660, A0=>nx26638, A1=>nx33670);
   ix17464 : mux21_ni port map ( Y=>nx17463, A0=>label_1_output(12), A1=>
      label_1_input_12, S0=>nx35609);
   ix6137 : mux21_ni port map ( Y=>nx6136, A0=>nx6132, A1=>
      label_1_input_state_machine_12, S0=>nx35957);
   ix17454 : mux21_ni port map ( Y=>nx17453, A0=>
      label_1_input_state_machine_12, A1=>mdr_data_out(12), S0=>nx35601);
   ix33676 : xnor2 port map ( Y=>nx33675, A0=>nx26636, A1=>nx33677);
   ix24334 : mux21_ni port map ( Y=>nx24333, A0=>nx13371, A1=>
      max_calc_ans1_14, S0=>nx35851);
   ix17207 : mux21_ni port map ( Y=>nx17206, A0=>max_calc_ans5_14, A1=>
      max_calc_ans6_14, S0=>nx35989);
   ix24344 : mux21_ni port map ( Y=>nx24343, A0=>max_calc_ans6_14, A1=>
      nx13371, S0=>nx36021);
   ix24354 : mux21_ni port map ( Y=>nx24353, A0=>max_calc_ans5_14, A1=>
      nx17196, S0=>nx35749);
   ix17197 : mux21 port map ( Y=>nx17196, A0=>nx27573, A1=>nx27763, S0=>
      nx35861);
   ix17257 : xor2 port map ( Y=>nx17256, A0=>nx33292, A1=>
      max_calc_comparator_first_inp1_14);
   ix33695 : xor2 port map ( Y=>nx33694, A0=>
      max_calc_comparator_first_inp2_13, A1=>
      max_calc_comparator_first_inp1_13);
   ix24474 : mux21_ni port map ( Y=>nx24473, A0=>
      max_calc_comparator_first_inp2_13, A1=>nx17370, S0=>nx36281);
   ix17371 : mux21_ni port map ( Y=>nx17370, A0=>nx17366, A1=>nx17278, S0=>
      nx35969);
   ix17279 : mux21_ni port map ( Y=>nx17278, A0=>max_calc_ans2_13, A1=>
      label_2_output(13), S0=>nx35989);
   ix24404 : mux21_ni port map ( Y=>nx24403, A0=>nx17268, A1=>
      max_calc_ans2_13, S0=>nx35851);
   ix17269 : mux21 port map ( Y=>nx17268, A0=>nx32869, A1=>nx32880, S0=>
      nx35899);
   ix17367 : mux21_ni port map ( Y=>nx17366, A0=>max_calc_ans8_13, A1=>
      max_calc_ans7_13, S0=>nx35989);
   ix24464 : mux21_ni port map ( Y=>nx24463, A0=>max_calc_ans7_13, A1=>
      nx17268, S0=>nx36021);
   ix24454 : mux21_ni port map ( Y=>nx24453, A0=>nx13375, A1=>
      max_calc_ans8_13, S0=>nx35869);
   ix17347 : mux21_ni port map ( Y=>nx13375, A0=>
      max_calc_comparator_first_inp2_13, A1=>
      max_calc_comparator_first_inp1_13, S0=>nx35905);
   ix24444 : mux21_ni port map ( Y=>nx24443, A0=>
      max_calc_comparator_first_inp1_13, A1=>nx17332, S0=>nx36281);
   ix17333 : mux21_ni port map ( Y=>nx17332, A0=>nx17328, A1=>nx17296, S0=>
      nx35969);
   ix17297 : mux21_ni port map ( Y=>nx17296, A0=>max_calc_ans1_13, A1=>
      label_1_output(13), S0=>nx35989);
   ix24414 : mux21_ni port map ( Y=>nx24413, A0=>nx13375, A1=>
      max_calc_ans1_13, S0=>nx35851);
   ix17329 : mux21_ni port map ( Y=>nx17328, A0=>max_calc_ans5_13, A1=>
      max_calc_ans6_13, S0=>nx35989);
   ix24424 : mux21_ni port map ( Y=>nx24423, A0=>max_calc_ans6_13, A1=>
      nx13375, S0=>nx36021);
   ix24434 : mux21_ni port map ( Y=>nx24433, A0=>max_calc_ans5_13, A1=>
      nx17318, S0=>nx35749);
   ix17319 : mux21 port map ( Y=>nx17318, A0=>nx27956, A1=>nx27960, S0=>
      nx35861);
   ix24554 : mux21_ni port map ( Y=>nx24553, A0=>
      max_calc_comparator_first_inp2_12, A1=>nx17492, S0=>nx36283);
   ix17493 : mux21_ni port map ( Y=>nx17492, A0=>nx17488, A1=>nx17400, S0=>
      nx35969);
   ix17401 : mux21_ni port map ( Y=>nx17400, A0=>max_calc_ans2_12, A1=>
      label_2_output(12), S0=>nx35989);
   ix24484 : mux21_ni port map ( Y=>nx24483, A0=>nx17390, A1=>
      max_calc_ans2_12, S0=>nx35851);
   ix17391 : mux21 port map ( Y=>nx17390, A0=>nx32894, A1=>nx32908, S0=>
      nx35899);
   ix17489 : mux21_ni port map ( Y=>nx17488, A0=>max_calc_ans8_12, A1=>
      max_calc_ans7_12, S0=>nx35991);
   ix24544 : mux21_ni port map ( Y=>nx24543, A0=>max_calc_ans7_12, A1=>
      nx17390, S0=>nx36021);
   ix24534 : mux21_ni port map ( Y=>nx24533, A0=>nx13376, A1=>
      max_calc_ans8_12, S0=>nx35869);
   ix17469 : mux21_ni port map ( Y=>nx13376, A0=>
      max_calc_comparator_first_inp2_12, A1=>
      max_calc_comparator_first_inp1_12, S0=>nx35905);
   ix24524 : mux21_ni port map ( Y=>nx24523, A0=>
      max_calc_comparator_first_inp1_12, A1=>nx17454, S0=>nx36283);
   ix17455 : mux21_ni port map ( Y=>nx17454, A0=>nx17450, A1=>nx17418, S0=>
      nx35969);
   ix17419 : mux21_ni port map ( Y=>nx17418, A0=>max_calc_ans1_12, A1=>
      label_1_output(12), S0=>nx35991);
   ix24494 : mux21_ni port map ( Y=>nx24493, A0=>nx13376, A1=>
      max_calc_ans1_12, S0=>nx35853);
   ix17451 : mux21_ni port map ( Y=>nx17450, A0=>max_calc_ans5_12, A1=>
      max_calc_ans6_12, S0=>nx35991);
   ix24504 : mux21_ni port map ( Y=>nx24503, A0=>max_calc_ans6_12, A1=>
      nx13376, S0=>nx36023);
   ix24514 : mux21_ni port map ( Y=>nx24513, A0=>max_calc_ans5_12, A1=>
      nx17440, S0=>nx35749);
   ix17441 : mux21 port map ( Y=>nx17440, A0=>nx27967, A1=>nx27974, S0=>
      nx35861);
   ix17501 : xor2 port map ( Y=>nx17500, A0=>nx33731, A1=>
      max_calc_comparator_first_inp1_12);
   ix33768 : xor2 port map ( Y=>nx33767, A0=>
      max_calc_comparator_first_inp2_11, A1=>
      max_calc_comparator_first_inp1_11);
   ix24634 : mux21_ni port map ( Y=>nx24633, A0=>
      max_calc_comparator_first_inp2_11, A1=>nx17614, S0=>nx36283);
   ix17615 : mux21_ni port map ( Y=>nx17614, A0=>nx17610, A1=>nx17522, S0=>
      nx35971);
   ix17523 : mux21_ni port map ( Y=>nx17522, A0=>max_calc_ans2_11, A1=>
      label_2_output(11), S0=>nx35991);
   ix24564 : mux21_ni port map ( Y=>nx24563, A0=>nx17512, A1=>
      max_calc_ans2_11, S0=>nx35853);
   ix17513 : mux21 port map ( Y=>nx17512, A0=>nx32925, A1=>nx32936, S0=>
      nx35899);
   ix17611 : mux21_ni port map ( Y=>nx17610, A0=>max_calc_ans8_11, A1=>
      max_calc_ans7_11, S0=>nx35991);
   ix24624 : mux21_ni port map ( Y=>nx24623, A0=>max_calc_ans7_11, A1=>
      nx17512, S0=>nx36023);
   ix24614 : mux21_ni port map ( Y=>nx24613, A0=>nx13377, A1=>
      max_calc_ans8_11, S0=>nx35869);
   ix17591 : mux21_ni port map ( Y=>nx13377, A0=>
      max_calc_comparator_first_inp2_11, A1=>
      max_calc_comparator_first_inp1_11, S0=>nx35905);
   ix24604 : mux21_ni port map ( Y=>nx24603, A0=>
      max_calc_comparator_first_inp1_11, A1=>nx17576, S0=>nx36283);
   ix17577 : mux21_ni port map ( Y=>nx17576, A0=>nx17572, A1=>nx17540, S0=>
      nx35971);
   ix17541 : mux21_ni port map ( Y=>nx17540, A0=>max_calc_ans1_11, A1=>
      label_1_output(11), S0=>nx35991);
   ix24574 : mux21_ni port map ( Y=>nx24573, A0=>nx13377, A1=>
      max_calc_ans1_11, S0=>nx35853);
   ix17573 : mux21_ni port map ( Y=>nx17572, A0=>max_calc_ans5_11, A1=>
      max_calc_ans6_11, S0=>nx35991);
   ix24584 : mux21_ni port map ( Y=>nx24583, A0=>max_calc_ans6_11, A1=>
      nx13377, S0=>nx36023);
   ix24594 : mux21_ni port map ( Y=>nx24593, A0=>max_calc_ans5_11, A1=>
      nx17562, S0=>nx35749);
   ix17563 : mux21 port map ( Y=>nx17562, A0=>nx27984, A1=>nx27988, S0=>
      nx35861);
   ix24714 : mux21_ni port map ( Y=>nx24713, A0=>
      max_calc_comparator_first_inp2_10, A1=>nx17736, S0=>nx36283);
   ix17737 : mux21_ni port map ( Y=>nx17736, A0=>nx17732, A1=>nx17644, S0=>
      nx35971);
   ix17645 : mux21_ni port map ( Y=>nx17644, A0=>max_calc_ans2_10, A1=>
      label_2_output(10), S0=>nx35993);
   ix24644 : mux21_ni port map ( Y=>nx24643, A0=>nx17634, A1=>
      max_calc_ans2_10, S0=>nx35853);
   ix17635 : mux21 port map ( Y=>nx17634, A0=>nx32950, A1=>nx32964, S0=>
      nx35899);
   ix17733 : mux21_ni port map ( Y=>nx17732, A0=>max_calc_ans8_10, A1=>
      max_calc_ans7_10, S0=>nx35993);
   ix24704 : mux21_ni port map ( Y=>nx24703, A0=>max_calc_ans7_10, A1=>
      nx17634, S0=>nx36023);
   ix24694 : mux21_ni port map ( Y=>nx24693, A0=>nx13379, A1=>
      max_calc_ans8_10, S0=>nx35869);
   ix17713 : mux21_ni port map ( Y=>nx13379, A0=>
      max_calc_comparator_first_inp2_10, A1=>
      max_calc_comparator_first_inp1_10, S0=>nx35905);
   ix24684 : mux21_ni port map ( Y=>nx24683, A0=>
      max_calc_comparator_first_inp1_10, A1=>nx17698, S0=>nx36283);
   ix17699 : mux21_ni port map ( Y=>nx17698, A0=>nx17694, A1=>nx17662, S0=>
      nx35971);
   ix17663 : mux21_ni port map ( Y=>nx17662, A0=>max_calc_ans1_10, A1=>
      label_1_output(10), S0=>nx35993);
   ix24654 : mux21_ni port map ( Y=>nx24653, A0=>nx13379, A1=>
      max_calc_ans1_10, S0=>nx35853);
   ix17695 : mux21_ni port map ( Y=>nx17694, A0=>max_calc_ans5_10, A1=>
      max_calc_ans6_10, S0=>nx35993);
   ix24664 : mux21_ni port map ( Y=>nx24663, A0=>max_calc_ans6_10, A1=>
      nx13379, S0=>nx36023);
   ix24674 : mux21_ni port map ( Y=>nx24673, A0=>max_calc_ans5_10, A1=>
      nx17684, S0=>nx35749);
   ix17685 : mux21 port map ( Y=>nx17684, A0=>nx27995, A1=>nx28002, S0=>
      nx35861);
   ix17745 : xor2 port map ( Y=>nx17744, A0=>nx33804, A1=>
      max_calc_comparator_first_inp1_10);
   ix33841 : xor2 port map ( Y=>nx33840, A0=>
      max_calc_comparator_first_inp2_9, A1=>max_calc_comparator_first_inp1_9
   );
   ix24794 : mux21_ni port map ( Y=>nx24793, A0=>
      max_calc_comparator_first_inp2_9, A1=>nx17858, S0=>nx36283);
   ix17859 : mux21_ni port map ( Y=>nx17858, A0=>nx17854, A1=>nx17766, S0=>
      nx35971);
   ix17767 : mux21_ni port map ( Y=>nx17766, A0=>max_calc_ans2_9, A1=>
      label_2_output(9), S0=>nx35993);
   ix24724 : mux21_ni port map ( Y=>nx24723, A0=>nx17756, A1=>
      max_calc_ans2_9, S0=>nx35853);
   ix17757 : mux21 port map ( Y=>nx17756, A0=>nx32981, A1=>nx32992, S0=>
      nx35899);
   ix17855 : mux21_ni port map ( Y=>nx17854, A0=>max_calc_ans8_9, A1=>
      max_calc_ans7_9, S0=>nx35993);
   ix24784 : mux21_ni port map ( Y=>nx24783, A0=>max_calc_ans7_9, A1=>
      nx17756, S0=>nx36023);
   ix24774 : mux21_ni port map ( Y=>nx24773, A0=>nx13381, A1=>
      max_calc_ans8_9, S0=>nx35871);
   ix17835 : mux21_ni port map ( Y=>nx13381, A0=>
      max_calc_comparator_first_inp2_9, A1=>max_calc_comparator_first_inp1_9, 
      S0=>nx35905);
   ix24764 : mux21_ni port map ( Y=>nx24763, A0=>
      max_calc_comparator_first_inp1_9, A1=>nx17820, S0=>nx36285);
   ix17821 : mux21_ni port map ( Y=>nx17820, A0=>nx17816, A1=>nx17784, S0=>
      nx35971);
   ix17785 : mux21_ni port map ( Y=>nx17784, A0=>max_calc_ans1_9, A1=>
      label_1_output(9), S0=>nx35993);
   ix24734 : mux21_ni port map ( Y=>nx24733, A0=>nx13381, A1=>
      max_calc_ans1_9, S0=>nx35853);
   ix17817 : mux21_ni port map ( Y=>nx17816, A0=>max_calc_ans5_9, A1=>
      max_calc_ans6_9, S0=>nx35995);
   ix24744 : mux21_ni port map ( Y=>nx24743, A0=>max_calc_ans6_9, A1=>
      nx13381, S0=>nx36023);
   ix24754 : mux21_ni port map ( Y=>nx24753, A0=>max_calc_ans5_9, A1=>
      nx17806, S0=>nx35749);
   ix17807 : mux21 port map ( Y=>nx17806, A0=>nx28012, A1=>nx28016, S0=>
      nx35861);
   ix24874 : mux21_ni port map ( Y=>nx24873, A0=>
      max_calc_comparator_first_inp2_8, A1=>nx17980, S0=>nx36285);
   ix17981 : mux21_ni port map ( Y=>nx17980, A0=>nx17976, A1=>nx17888, S0=>
      nx35971);
   ix17889 : mux21_ni port map ( Y=>nx17888, A0=>max_calc_ans2_8, A1=>
      label_2_output(8), S0=>nx35995);
   ix24804 : mux21_ni port map ( Y=>nx24803, A0=>nx17878, A1=>
      max_calc_ans2_8, S0=>nx35855);
   ix17879 : mux21 port map ( Y=>nx17878, A0=>nx33006, A1=>nx33020, S0=>
      nx35901);
   ix17977 : mux21_ni port map ( Y=>nx17976, A0=>max_calc_ans8_8, A1=>
      max_calc_ans7_8, S0=>nx35995);
   ix24864 : mux21_ni port map ( Y=>nx24863, A0=>max_calc_ans7_8, A1=>
      nx17878, S0=>nx36025);
   ix24854 : mux21_ni port map ( Y=>nx24853, A0=>nx13383, A1=>
      max_calc_ans8_8, S0=>nx35871);
   ix17957 : mux21_ni port map ( Y=>nx13383, A0=>
      max_calc_comparator_first_inp2_8, A1=>max_calc_comparator_first_inp1_8, 
      S0=>nx35907);
   ix24844 : mux21_ni port map ( Y=>nx24843, A0=>
      max_calc_comparator_first_inp1_8, A1=>nx17942, S0=>nx36285);
   ix17943 : mux21_ni port map ( Y=>nx17942, A0=>nx17938, A1=>nx17906, S0=>
      nx35973);
   ix17907 : mux21_ni port map ( Y=>nx17906, A0=>max_calc_ans1_8, A1=>
      label_1_output(8), S0=>nx35995);
   ix24814 : mux21_ni port map ( Y=>nx24813, A0=>nx13383, A1=>
      max_calc_ans1_8, S0=>nx35855);
   ix17939 : mux21_ni port map ( Y=>nx17938, A0=>max_calc_ans5_8, A1=>
      max_calc_ans6_8, S0=>nx35995);
   ix24824 : mux21_ni port map ( Y=>nx24823, A0=>max_calc_ans6_8, A1=>
      nx13383, S0=>nx36025);
   ix24834 : mux21_ni port map ( Y=>nx24833, A0=>max_calc_ans5_8, A1=>
      nx17928, S0=>nx35751);
   ix17929 : mux21 port map ( Y=>nx17928, A0=>nx28023, A1=>nx28030, S0=>
      nx35863);
   ix17989 : xor2 port map ( Y=>nx17988, A0=>nx33877, A1=>
      max_calc_comparator_first_inp1_8);
   ix33914 : xor2 port map ( Y=>nx33913, A0=>
      max_calc_comparator_first_inp2_7, A1=>max_calc_comparator_first_inp1_7
   );
   ix24954 : mux21_ni port map ( Y=>nx24953, A0=>
      max_calc_comparator_first_inp2_7, A1=>nx18102, S0=>nx36285);
   ix18103 : mux21_ni port map ( Y=>nx18102, A0=>nx18098, A1=>nx18010, S0=>
      nx35973);
   ix18011 : mux21_ni port map ( Y=>nx18010, A0=>max_calc_ans2_7, A1=>
      label_2_output(7), S0=>nx35995);
   ix24884 : mux21_ni port map ( Y=>nx24883, A0=>nx18000, A1=>
      max_calc_ans2_7, S0=>nx35855);
   ix18001 : mux21 port map ( Y=>nx18000, A0=>nx33037, A1=>nx33048, S0=>
      nx35901);
   ix18099 : mux21_ni port map ( Y=>nx18098, A0=>max_calc_ans8_7, A1=>
      max_calc_ans7_7, S0=>nx35995);
   ix24944 : mux21_ni port map ( Y=>nx24943, A0=>max_calc_ans7_7, A1=>
      nx18000, S0=>nx36025);
   ix24934 : mux21_ni port map ( Y=>nx24933, A0=>nx13385, A1=>
      max_calc_ans8_7, S0=>nx35871);
   ix18079 : mux21_ni port map ( Y=>nx13385, A0=>
      max_calc_comparator_first_inp2_7, A1=>max_calc_comparator_first_inp1_7, 
      S0=>nx35907);
   ix24924 : mux21_ni port map ( Y=>nx24923, A0=>
      max_calc_comparator_first_inp1_7, A1=>nx18064, S0=>nx36285);
   ix18065 : mux21_ni port map ( Y=>nx18064, A0=>nx18060, A1=>nx18028, S0=>
      nx35973);
   ix18029 : mux21_ni port map ( Y=>nx18028, A0=>max_calc_ans1_7, A1=>
      label_1_output(7), S0=>nx35997);
   ix24894 : mux21_ni port map ( Y=>nx24893, A0=>nx13385, A1=>
      max_calc_ans1_7, S0=>nx35855);
   ix18061 : mux21_ni port map ( Y=>nx18060, A0=>max_calc_ans5_7, A1=>
      max_calc_ans6_7, S0=>nx35997);
   ix24904 : mux21_ni port map ( Y=>nx24903, A0=>max_calc_ans6_7, A1=>
      nx13385, S0=>nx36025);
   ix24914 : mux21_ni port map ( Y=>nx24913, A0=>max_calc_ans5_7, A1=>
      nx18050, S0=>nx35751);
   ix18051 : mux21 port map ( Y=>nx18050, A0=>nx28040, A1=>nx28044, S0=>
      nx35863);
   ix25034 : mux21_ni port map ( Y=>nx25033, A0=>
      max_calc_comparator_first_inp2_6, A1=>nx18224, S0=>nx36285);
   ix18225 : mux21_ni port map ( Y=>nx18224, A0=>nx18220, A1=>nx18132, S0=>
      nx35973);
   ix18133 : mux21_ni port map ( Y=>nx18132, A0=>max_calc_ans2_6, A1=>
      label_2_output(6), S0=>nx35997);
   ix24964 : mux21_ni port map ( Y=>nx24963, A0=>nx18122, A1=>
      max_calc_ans2_6, S0=>nx35855);
   ix18123 : mux21 port map ( Y=>nx18122, A0=>nx33062, A1=>nx33076, S0=>
      nx35901);
   ix18221 : mux21_ni port map ( Y=>nx18220, A0=>max_calc_ans8_6, A1=>
      max_calc_ans7_6, S0=>nx35997);
   ix25024 : mux21_ni port map ( Y=>nx25023, A0=>max_calc_ans7_6, A1=>
      nx18122, S0=>nx36025);
   ix25014 : mux21_ni port map ( Y=>nx25013, A0=>nx13386, A1=>
      max_calc_ans8_6, S0=>nx35871);
   ix18201 : mux21_ni port map ( Y=>nx13386, A0=>
      max_calc_comparator_first_inp2_6, A1=>max_calc_comparator_first_inp1_6, 
      S0=>nx35907);
   ix25004 : mux21_ni port map ( Y=>nx25003, A0=>
      max_calc_comparator_first_inp1_6, A1=>nx18186, S0=>nx36285);
   ix18187 : mux21_ni port map ( Y=>nx18186, A0=>nx18182, A1=>nx18150, S0=>
      nx35973);
   ix18151 : mux21_ni port map ( Y=>nx18150, A0=>max_calc_ans1_6, A1=>
      label_1_output(6), S0=>nx35997);
   ix24974 : mux21_ni port map ( Y=>nx24973, A0=>nx13386, A1=>
      max_calc_ans1_6, S0=>nx35855);
   ix18183 : mux21_ni port map ( Y=>nx18182, A0=>max_calc_ans5_6, A1=>
      max_calc_ans6_6, S0=>nx35997);
   ix24984 : mux21_ni port map ( Y=>nx24983, A0=>max_calc_ans6_6, A1=>
      nx13386, S0=>nx36025);
   ix24994 : mux21_ni port map ( Y=>nx24993, A0=>max_calc_ans5_6, A1=>
      nx18172, S0=>nx35751);
   ix18173 : mux21 port map ( Y=>nx18172, A0=>nx28051, A1=>nx28058, S0=>
      nx35863);
   ix18233 : xor2 port map ( Y=>nx18232, A0=>nx33950, A1=>
      max_calc_comparator_first_inp1_6);
   ix33987 : xor2 port map ( Y=>nx33986, A0=>
      max_calc_comparator_first_inp2_5, A1=>max_calc_comparator_first_inp1_5
   );
   ix25114 : mux21_ni port map ( Y=>nx25113, A0=>
      max_calc_comparator_first_inp2_5, A1=>nx18346, S0=>nx36287);
   ix18347 : mux21_ni port map ( Y=>nx18346, A0=>nx18342, A1=>nx18254, S0=>
      nx35973);
   ix18255 : mux21_ni port map ( Y=>nx18254, A0=>max_calc_ans2_5, A1=>
      label_2_output(5), S0=>nx35997);
   ix25044 : mux21_ni port map ( Y=>nx25043, A0=>nx18244, A1=>
      max_calc_ans2_5, S0=>nx35855);
   ix18245 : mux21 port map ( Y=>nx18244, A0=>nx33093, A1=>nx33104, S0=>
      nx35901);
   ix18343 : mux21_ni port map ( Y=>nx18342, A0=>max_calc_ans8_5, A1=>
      max_calc_ans7_5, S0=>nx35189);
   ix25104 : mux21_ni port map ( Y=>nx25103, A0=>max_calc_ans7_5, A1=>
      nx18244, S0=>nx36025);
   ix25094 : mux21_ni port map ( Y=>nx25093, A0=>nx13387, A1=>
      max_calc_ans8_5, S0=>nx35871);
   ix18323 : mux21_ni port map ( Y=>nx13387, A0=>
      max_calc_comparator_first_inp2_5, A1=>max_calc_comparator_first_inp1_5, 
      S0=>nx35907);
   ix25084 : mux21_ni port map ( Y=>nx25083, A0=>
      max_calc_comparator_first_inp1_5, A1=>nx18308, S0=>nx36287);
   ix18309 : mux21_ni port map ( Y=>nx18308, A0=>nx18304, A1=>nx18272, S0=>
      nx35973);
   ix18273 : mux21_ni port map ( Y=>nx18272, A0=>max_calc_ans1_5, A1=>
      label_1_output(5), S0=>nx35189);
   ix25054 : mux21_ni port map ( Y=>nx25053, A0=>nx13387, A1=>
      max_calc_ans1_5, S0=>nx35857);
   ix18305 : mux21_ni port map ( Y=>nx18304, A0=>max_calc_ans5_5, A1=>
      max_calc_ans6_5, S0=>nx35189);
   ix25064 : mux21_ni port map ( Y=>nx25063, A0=>max_calc_ans6_5, A1=>
      nx13387, S0=>nx36027);
   ix25074 : mux21_ni port map ( Y=>nx25073, A0=>max_calc_ans5_5, A1=>
      nx18294, S0=>nx35751);
   ix18295 : mux21 port map ( Y=>nx18294, A0=>nx28068, A1=>nx28072, S0=>
      nx35863);
   ix25194 : mux21_ni port map ( Y=>nx25193, A0=>
      max_calc_comparator_first_inp2_4, A1=>nx18468, S0=>nx36287);
   ix18469 : mux21_ni port map ( Y=>nx18468, A0=>nx18464, A1=>nx18376, S0=>
      nx35975);
   ix18377 : mux21_ni port map ( Y=>nx18376, A0=>max_calc_ans2_4, A1=>
      label_2_output(4), S0=>nx35189);
   ix25124 : mux21_ni port map ( Y=>nx25123, A0=>nx18366, A1=>
      max_calc_ans2_4, S0=>nx35857);
   ix18367 : mux21 port map ( Y=>nx18366, A0=>nx33118, A1=>nx33132, S0=>
      nx35901);
   ix18465 : mux21_ni port map ( Y=>nx18464, A0=>max_calc_ans8_4, A1=>
      max_calc_ans7_4, S0=>nx35189);
   ix25184 : mux21_ni port map ( Y=>nx25183, A0=>max_calc_ans7_4, A1=>
      nx18366, S0=>nx36027);
   ix25174 : mux21_ni port map ( Y=>nx25173, A0=>nx13388, A1=>
      max_calc_ans8_4, S0=>nx35871);
   ix18445 : mux21_ni port map ( Y=>nx13388, A0=>
      max_calc_comparator_first_inp2_4, A1=>max_calc_comparator_first_inp1_4, 
      S0=>nx35907);
   ix25164 : mux21_ni port map ( Y=>nx25163, A0=>
      max_calc_comparator_first_inp1_4, A1=>nx18430, S0=>nx36287);
   ix18431 : mux21_ni port map ( Y=>nx18430, A0=>nx18426, A1=>nx18394, S0=>
      nx35975);
   ix18395 : mux21_ni port map ( Y=>nx18394, A0=>max_calc_ans1_4, A1=>
      label_1_output(4), S0=>nx35189);
   ix25134 : mux21_ni port map ( Y=>nx25133, A0=>nx13388, A1=>
      max_calc_ans1_4, S0=>nx35857);
   ix18427 : mux21_ni port map ( Y=>nx18426, A0=>max_calc_ans5_4, A1=>
      max_calc_ans6_4, S0=>nx35189);
   ix25144 : mux21_ni port map ( Y=>nx25143, A0=>max_calc_ans6_4, A1=>
      nx13388, S0=>nx36027);
   ix25154 : mux21_ni port map ( Y=>nx25153, A0=>max_calc_ans5_4, A1=>
      nx18416, S0=>nx35751);
   ix18417 : mux21 port map ( Y=>nx18416, A0=>nx28079, A1=>nx28086, S0=>
      nx35863);
   ix18477 : xor2 port map ( Y=>nx18476, A0=>nx34023, A1=>
      max_calc_comparator_first_inp1_4);
   ix34060 : xor2 port map ( Y=>nx34059, A0=>
      max_calc_comparator_first_inp2_3, A1=>max_calc_comparator_first_inp1_3
   );
   ix25274 : mux21_ni port map ( Y=>nx25273, A0=>
      max_calc_comparator_first_inp2_3, A1=>nx18590, S0=>nx36287);
   ix18591 : mux21_ni port map ( Y=>nx18590, A0=>nx18586, A1=>nx18498, S0=>
      nx35975);
   ix18499 : mux21_ni port map ( Y=>nx18498, A0=>max_calc_ans2_3, A1=>
      label_2_output(3), S0=>nx35999);
   ix25204 : mux21_ni port map ( Y=>nx25203, A0=>nx18488, A1=>
      max_calc_ans2_3, S0=>nx35857);
   ix18489 : mux21 port map ( Y=>nx18488, A0=>nx33149, A1=>nx33160, S0=>
      nx35901);
   ix18587 : mux21_ni port map ( Y=>nx18586, A0=>max_calc_ans8_3, A1=>
      max_calc_ans7_3, S0=>nx35999);
   ix25264 : mux21_ni port map ( Y=>nx25263, A0=>max_calc_ans7_3, A1=>
      nx18488, S0=>nx36027);
   ix25254 : mux21_ni port map ( Y=>nx25253, A0=>nx13389, A1=>
      max_calc_ans8_3, S0=>nx35871);
   ix18567 : mux21_ni port map ( Y=>nx13389, A0=>
      max_calc_comparator_first_inp2_3, A1=>max_calc_comparator_first_inp1_3, 
      S0=>nx35907);
   ix25244 : mux21_ni port map ( Y=>nx25243, A0=>
      max_calc_comparator_first_inp1_3, A1=>nx18552, S0=>nx36287);
   ix18553 : mux21_ni port map ( Y=>nx18552, A0=>nx18548, A1=>nx18516, S0=>
      nx35975);
   ix18517 : mux21_ni port map ( Y=>nx18516, A0=>max_calc_ans1_3, A1=>
      label_1_output(3), S0=>nx35999);
   ix25214 : mux21_ni port map ( Y=>nx25213, A0=>nx13389, A1=>
      max_calc_ans1_3, S0=>nx35857);
   ix18549 : mux21_ni port map ( Y=>nx18548, A0=>max_calc_ans5_3, A1=>
      max_calc_ans6_3, S0=>nx35999);
   ix25224 : mux21_ni port map ( Y=>nx25223, A0=>max_calc_ans6_3, A1=>
      nx13389, S0=>nx36027);
   ix25234 : mux21_ni port map ( Y=>nx25233, A0=>max_calc_ans5_3, A1=>
      nx18538, S0=>nx35751);
   ix18539 : mux21 port map ( Y=>nx18538, A0=>nx28096, A1=>nx28100, S0=>
      nx35863);
   ix25354 : mux21_ni port map ( Y=>nx25353, A0=>
      max_calc_comparator_first_inp2_2, A1=>nx18712, S0=>nx36287);
   ix18713 : mux21_ni port map ( Y=>nx18712, A0=>nx18708, A1=>nx18620, S0=>
      nx35975);
   ix18621 : mux21_ni port map ( Y=>nx18620, A0=>max_calc_ans2_2, A1=>
      label_2_output(2), S0=>nx35999);
   ix25284 : mux21_ni port map ( Y=>nx25283, A0=>nx18610, A1=>
      max_calc_ans2_2, S0=>nx35857);
   ix18611 : mux21 port map ( Y=>nx18610, A0=>nx33174, A1=>nx33188, S0=>
      nx35901);
   ix18709 : mux21_ni port map ( Y=>nx18708, A0=>max_calc_ans8_2, A1=>
      max_calc_ans7_2, S0=>nx35999);
   ix25344 : mux21_ni port map ( Y=>nx25343, A0=>max_calc_ans7_2, A1=>
      nx18610, S0=>nx36027);
   ix25334 : mux21_ni port map ( Y=>nx25333, A0=>nx13391, A1=>
      max_calc_ans8_2, S0=>nx35873);
   ix18689 : mux21_ni port map ( Y=>nx13391, A0=>
      max_calc_comparator_first_inp2_2, A1=>max_calc_comparator_first_inp1_2, 
      S0=>nx35907);
   ix25324 : mux21_ni port map ( Y=>nx25323, A0=>
      max_calc_comparator_first_inp1_2, A1=>nx18674, S0=>nx36289);
   ix18675 : mux21_ni port map ( Y=>nx18674, A0=>nx18670, A1=>nx18638, S0=>
      nx35975);
   ix18639 : mux21_ni port map ( Y=>nx18638, A0=>max_calc_ans1_2, A1=>
      label_1_output(2), S0=>nx35999);
   ix25294 : mux21_ni port map ( Y=>nx25293, A0=>nx13391, A1=>
      max_calc_ans1_2, S0=>nx35857);
   ix18671 : mux21_ni port map ( Y=>nx18670, A0=>max_calc_ans5_2, A1=>
      max_calc_ans6_2, S0=>nx36001);
   ix25304 : mux21_ni port map ( Y=>nx25303, A0=>max_calc_ans6_2, A1=>
      nx13391, S0=>nx36027);
   ix25314 : mux21_ni port map ( Y=>nx25313, A0=>max_calc_ans5_2, A1=>
      nx18660, S0=>nx35751);
   ix18661 : mux21 port map ( Y=>nx18660, A0=>nx28107, A1=>nx28114, S0=>
      nx35863);
   ix18721 : xor2 port map ( Y=>nx18720, A0=>nx34096, A1=>
      max_calc_comparator_first_inp1_2);
   ix25434 : mux21_ni port map ( Y=>nx25433, A0=>
      max_calc_comparator_first_inp2_1, A1=>nx18834, S0=>nx36289);
   ix18835 : mux21_ni port map ( Y=>nx18834, A0=>nx18830, A1=>nx18742, S0=>
      nx35975);
   ix18743 : mux21_ni port map ( Y=>nx18742, A0=>max_calc_ans2_1, A1=>
      label_2_output(1), S0=>nx36001);
   ix25364 : mux21_ni port map ( Y=>nx25363, A0=>nx18732, A1=>
      max_calc_ans2_1, S0=>nx35859);
   ix18733 : mux21 port map ( Y=>nx18732, A0=>nx33203, A1=>nx33214, S0=>
      nx35903);
   ix18831 : mux21_ni port map ( Y=>nx18830, A0=>max_calc_ans8_1, A1=>
      max_calc_ans7_1, S0=>nx36001);
   ix25424 : mux21_ni port map ( Y=>nx25423, A0=>max_calc_ans7_1, A1=>
      nx18732, S0=>nx36029);
   ix25414 : mux21_ni port map ( Y=>nx25413, A0=>nx13393, A1=>
      max_calc_ans8_1, S0=>nx35873);
   ix18811 : mux21_ni port map ( Y=>nx13393, A0=>
      max_calc_comparator_first_inp2_1, A1=>max_calc_comparator_first_inp1_1, 
      S0=>nx35909);
   ix25404 : mux21_ni port map ( Y=>nx25403, A0=>
      max_calc_comparator_first_inp1_1, A1=>nx18796, S0=>nx36289);
   ix18797 : mux21_ni port map ( Y=>nx18796, A0=>nx18792, A1=>nx18760, S0=>
      nx35185);
   ix18761 : mux21_ni port map ( Y=>nx18760, A0=>max_calc_ans1_1, A1=>
      label_1_output(1), S0=>nx36001);
   ix25374 : mux21_ni port map ( Y=>nx25373, A0=>nx13393, A1=>
      max_calc_ans1_1, S0=>nx35859);
   ix18793 : mux21_ni port map ( Y=>nx18792, A0=>max_calc_ans5_1, A1=>
      max_calc_ans6_1, S0=>nx36001);
   ix25384 : mux21_ni port map ( Y=>nx25383, A0=>max_calc_ans6_1, A1=>
      nx13393, S0=>nx36029);
   ix25394 : mux21_ni port map ( Y=>nx25393, A0=>max_calc_ans5_1, A1=>
      nx18782, S0=>nx35753);
   ix18783 : mux21 port map ( Y=>nx18782, A0=>nx28122, A1=>nx28126, S0=>
      nx35865);
   ix18843 : xor2 port map ( Y=>nx18842, A0=>
      max_calc_comparator_first_inp2_1, A1=>nx34162);
   ix25554 : mux21_ni port map ( Y=>nx25553, A0=>
      max_calc_comparator_first_inp2_15, A1=>nx19132, S0=>nx36289);
   ix19133 : mux21_ni port map ( Y=>nx19132, A0=>nx19128, A1=>nx19040, S0=>
      nx35185);
   ix19041 : mux21_ni port map ( Y=>nx19040, A0=>max_calc_ans2_15, A1=>
      label_2_output(15), S0=>nx36001);
   ix16664 : mux21_ni port map ( Y=>nx16663, A0=>label_2_output(15), A1=>
      label_2_input_15, S0=>nx35609);
   ix4889 : mux21_ni port map ( Y=>nx4888, A0=>nx4884, A1=>
      label_2_input_state_machine_15, S0=>nx35171);
   ix15824 : mux21_ni port map ( Y=>nx15823, A0=>
      label_2_input_state_machine_15, A1=>mdr_data_out(31), S0=>nx35601);
   ix34183 : xor2 port map ( Y=>nx34182, A0=>nx28594, A1=>label_2_output(15)
   );
   ix25484 : mux21_ni port map ( Y=>nx25483, A0=>nx19030, A1=>
      max_calc_ans2_15, S0=>nx35859);
   ix19031 : mux21 port map ( Y=>nx19030, A0=>nx33232, A1=>nx33257, S0=>
      nx35903);
   ix19129 : mux21_ni port map ( Y=>nx19128, A0=>max_calc_ans8_15, A1=>
      max_calc_ans7_15, S0=>nx36001);
   ix25544 : mux21_ni port map ( Y=>nx25543, A0=>max_calc_ans7_15, A1=>
      nx19030, S0=>nx36029);
   ix25534 : mux21_ni port map ( Y=>nx25533, A0=>nx13395, A1=>
      max_calc_ans8_15, S0=>nx35873);
   ix19109 : mux21_ni port map ( Y=>nx13395, A0=>
      max_calc_comparator_first_inp2_15, A1=>
      max_calc_comparator_first_inp1_15, S0=>nx35909);
   ix25524 : mux21_ni port map ( Y=>nx25523, A0=>
      max_calc_comparator_first_inp1_15, A1=>nx19094, S0=>nx36289);
   ix19095 : mux21_ni port map ( Y=>nx19094, A0=>nx19090, A1=>nx19058, S0=>
      nx35185);
   ix19059 : mux21_ni port map ( Y=>nx19058, A0=>max_calc_ans1_15, A1=>
      label_1_output(15), S0=>nx35191);
   ix17514 : mux21_ni port map ( Y=>nx17513, A0=>label_1_output(15), A1=>
      label_1_input_15, S0=>nx35609);
   ix6227 : mux21_ni port map ( Y=>nx6226, A0=>nx6222, A1=>
      label_1_input_state_machine_15, S0=>nx35171);
   ix16674 : mux21_ni port map ( Y=>nx16673, A0=>
      label_1_input_state_machine_15, A1=>mdr_data_out(15), S0=>nx35601);
   ix34210 : xor2 port map ( Y=>nx34209, A0=>nx26634, A1=>label_1_output(15)
   );
   ix25494 : mux21_ni port map ( Y=>nx25493, A0=>nx13395, A1=>
      max_calc_ans1_15, S0=>nx35859);
   ix19091 : mux21_ni port map ( Y=>nx19090, A0=>max_calc_ans5_15, A1=>
      max_calc_ans6_15, S0=>nx35191);
   ix25504 : mux21_ni port map ( Y=>nx25503, A0=>max_calc_ans6_15, A1=>
      nx13395, S0=>nx36029);
   ix25514 : mux21_ni port map ( Y=>nx25513, A0=>max_calc_ans5_15, A1=>
      nx19080, S0=>nx35753);
   ix19081 : mux21 port map ( Y=>nx19080, A0=>nx28137, A1=>nx28155, S0=>
      nx35865);
   ix34227 : nor04 port map ( Y=>nx6342, A0=>nx35737, A1=>nx26180, A2=>
      nx26203, A3=>nx35711);
   ix6341 : nand02 port map ( Y=>nx35711, A0=>nx35191, A1=>nx26188);
   ix25574 : mux21_ni port map ( Y=>nx25573, A0=>answer_1_EXMPLR, A1=>
      nx13393, S0=>nx35741);
   ix25584 : mux21_ni port map ( Y=>nx25583, A0=>answer_2_EXMPLR, A1=>
      nx13391, S0=>nx35741);
   ix25594 : mux21_ni port map ( Y=>nx25593, A0=>answer_3_EXMPLR, A1=>
      nx13389, S0=>nx35741);
   ix25604 : mux21_ni port map ( Y=>nx25603, A0=>answer_4_EXMPLR, A1=>
      nx13388, S0=>nx35741);
   ix25614 : mux21_ni port map ( Y=>nx25613, A0=>answer_5_EXMPLR, A1=>
      nx13387, S0=>nx35741);
   ix25624 : mux21_ni port map ( Y=>nx25623, A0=>answer_6_EXMPLR, A1=>
      nx13386, S0=>nx35743);
   ix25634 : mux21_ni port map ( Y=>nx25633, A0=>answer_7_EXMPLR, A1=>
      nx13385, S0=>nx35743);
   ix25644 : mux21_ni port map ( Y=>nx25643, A0=>answer_8_EXMPLR, A1=>
      nx13383, S0=>nx35743);
   ix25654 : mux21_ni port map ( Y=>nx25653, A0=>answer_9_EXMPLR, A1=>
      nx13381, S0=>nx35743);
   ix25664 : mux21_ni port map ( Y=>nx25663, A0=>answer_10_EXMPLR, A1=>
      nx13379, S0=>nx35743);
   ix25674 : mux21_ni port map ( Y=>nx25673, A0=>answer_11_EXMPLR, A1=>
      nx13377, S0=>nx35743);
   ix25684 : mux21_ni port map ( Y=>nx25683, A0=>answer_12_EXMPLR, A1=>
      nx13376, S0=>nx35743);
   ix25694 : mux21_ni port map ( Y=>nx25693, A0=>answer_13_EXMPLR, A1=>
      nx13375, S0=>nx35745);
   ix25704 : mux21_ni port map ( Y=>nx25703, A0=>answer_14_EXMPLR, A1=>
      nx13371, S0=>nx35745);
   ix25714 : mux21_ni port map ( Y=>nx25713, A0=>answer_15_EXMPLR, A1=>
      nx13395, S0=>nx35745);
   ix191 : and02 port map ( Y=>nx190, A0=>nx12893, A1=>nx25907);
   ix19277 : nor02ii port map ( Y=>nx19276, A0=>nx38, A1=>nx12887);
   ix19241 : nor02ii port map ( Y=>nx19240, A0=>nx34380, A1=>nx26129);
   ix34381 : nor02ii port map ( Y=>nx34380, A0=>nx19232, A1=>nx12879);
   ix34584 : and02 port map ( Y=>nx34585, A0=>nx30681, A1=>nx35721);
   ix34586 : and02 port map ( Y=>nx34587, A0=>nx30681, A1=>nx35721);
   ix34616 : and02 port map ( Y=>nx34617, A0=>nx28752, A1=>nx35725);
   ix34618 : and02 port map ( Y=>nx34619, A0=>nx28752, A1=>nx35725);
   ix34648 : and02 port map ( Y=>nx34649, A0=>nx28309, A1=>nx35729);
   ix34650 : and02 port map ( Y=>nx34651, A0=>nx28309, A1=>nx35729);
   ix34680 : and02 port map ( Y=>nx34681, A0=>nx26349, A1=>nx35733);
   ix34682 : and02 port map ( Y=>nx34683, A0=>nx26349, A1=>nx35733);
   ix34860 : and02 port map ( Y=>nx34861, A0=>nx26828, A1=>nx35757);
   ix34862 : and02 port map ( Y=>nx34863, A0=>nx26828, A1=>nx35757);
   ix34892 : and02 port map ( Y=>nx34893, A0=>nx27267, A1=>nx35761);
   ix34894 : and02 port map ( Y=>nx34895, A0=>nx27267, A1=>nx35761);
   ix34952 : and02 port map ( Y=>nx34953, A0=>nx29195, A1=>nx35765);
   ix34954 : and02 port map ( Y=>nx34955, A0=>nx29195, A1=>nx35765);
   ix34984 : and02 port map ( Y=>nx34985, A0=>nx29636, A1=>nx35769);
   ix34986 : and02 port map ( Y=>nx34987, A0=>nx29636, A1=>nx35769);
   ix35024 : and02 port map ( Y=>nx35025, A0=>nx31124, A1=>nx35773);
   ix35026 : and02 port map ( Y=>nx35027, A0=>nx31124, A1=>nx35773);
   ix35056 : and02 port map ( Y=>nx35057, A0=>nx31563, A1=>nx35777);
   ix35058 : and02 port map ( Y=>nx35059, A0=>nx31563, A1=>nx35777);
   ix35712 : inv02 port map ( Y=>nx35713, A=>nx35149);
   ix35714 : inv02 port map ( Y=>nx35715, A=>nx35149);
   ix35716 : inv02 port map ( Y=>nx35717, A=>nx35149);
   ix35718 : inv01 port map ( Y=>nx35719, A=>nx30685);
   ix35720 : inv01 port map ( Y=>nx35721, A=>nx30685);
   ix35722 : inv01 port map ( Y=>nx35723, A=>nx28756);
   ix35724 : inv01 port map ( Y=>nx35725, A=>nx28756);
   ix35726 : inv01 port map ( Y=>nx35727, A=>nx28313);
   ix35728 : inv01 port map ( Y=>nx35729, A=>nx28313);
   ix35730 : inv01 port map ( Y=>nx35731, A=>nx26353);
   ix35732 : inv01 port map ( Y=>nx35733, A=>nx26353);
   ix35734 : inv02 port map ( Y=>nx35735, A=>nx36389);
   ix35736 : inv02 port map ( Y=>nx35737, A=>nx36389);
   ix35738 : inv01 port map ( Y=>nx35739, A=>nx6342);
   ix35740 : inv02 port map ( Y=>nx35741, A=>nx35739);
   ix35742 : inv02 port map ( Y=>nx35743, A=>nx35739);
   ix35744 : inv02 port map ( Y=>nx35745, A=>nx35739);
   ix35746 : inv02 port map ( Y=>nx35747, A=>nx26675);
   ix35748 : inv02 port map ( Y=>nx35749, A=>nx36381);
   ix35750 : inv02 port map ( Y=>nx35751, A=>nx36381);
   ix35752 : inv02 port map ( Y=>nx35753, A=>nx36381);
   ix35754 : inv01 port map ( Y=>nx35755, A=>nx26832);
   ix35756 : inv01 port map ( Y=>nx35757, A=>nx26832);
   ix35758 : inv01 port map ( Y=>nx35759, A=>nx27271);
   ix35760 : inv01 port map ( Y=>nx35761, A=>nx27271);
   ix35762 : inv01 port map ( Y=>nx35763, A=>nx29199);
   ix35764 : inv01 port map ( Y=>nx35765, A=>nx29199);
   ix35766 : inv01 port map ( Y=>nx35767, A=>nx29640);
   ix35768 : inv01 port map ( Y=>nx35769, A=>nx29640);
   ix35770 : inv01 port map ( Y=>nx35771, A=>nx31128);
   ix35772 : inv01 port map ( Y=>nx35773, A=>nx31128);
   ix35774 : inv01 port map ( Y=>nx35775, A=>nx31567);
   ix35776 : inv01 port map ( Y=>nx35777, A=>nx31567);
   ix35778 : inv02 port map ( Y=>nx35779, A=>state(1));
   ix35780 : inv02 port map ( Y=>nx35781, A=>state(1));
   ix35782 : inv02 port map ( Y=>nx35783, A=>state(2));
   ix35784 : inv02 port map ( Y=>nx35785, A=>state(2));
   ix35786 : buf02 port map ( Y=>nx35787, A=>nx25874);
   ix35788 : buf02 port map ( Y=>nx35789, A=>nx25874);
   ix35790 : inv01 port map ( Y=>nx35791, A=>sub_state(2));
   ix35792 : inv01 port map ( Y=>nx35793, A=>sub_state(2));
   ix35794 : buf02 port map ( Y=>nx35795, A=>nx25949);
   ix35796 : buf02 port map ( Y=>nx35797, A=>nx25949);
   ix35798 : inv02 port map ( Y=>nx35799, A=>nx34499);
   ix35800 : inv02 port map ( Y=>nx35801, A=>nx34499);
   ix35802 : buf02 port map ( Y=>nx35803, A=>nx26323);
   ix35804 : buf02 port map ( Y=>nx35805, A=>nx26323);
   ix35806 : buf02 port map ( Y=>nx35807, A=>nx26802);
   ix35808 : buf02 port map ( Y=>nx35809, A=>nx26802);
   ix35810 : buf02 port map ( Y=>nx35811, A=>nx27241);
   ix35812 : buf02 port map ( Y=>nx35813, A=>nx27241);
   ix35814 : buf02 port map ( Y=>nx35815, A=>nx28283);
   ix35816 : buf02 port map ( Y=>nx35817, A=>nx28283);
   ix35818 : buf02 port map ( Y=>nx35819, A=>nx28726);
   ix35820 : buf02 port map ( Y=>nx35821, A=>nx28726);
   ix35822 : buf02 port map ( Y=>nx35823, A=>nx29169);
   ix35824 : buf02 port map ( Y=>nx35825, A=>nx29169);
   ix35826 : buf02 port map ( Y=>nx35827, A=>nx29610);
   ix35828 : buf02 port map ( Y=>nx35829, A=>nx29610);
   ix35830 : buf02 port map ( Y=>nx35831, A=>nx30655);
   ix35832 : buf02 port map ( Y=>nx35833, A=>nx30655);
   ix35834 : buf02 port map ( Y=>nx35835, A=>nx31098);
   ix35836 : buf02 port map ( Y=>nx35837, A=>nx31098);
   ix35838 : buf02 port map ( Y=>nx35839, A=>nx31537);
   ix35840 : buf02 port map ( Y=>nx35841, A=>nx31537);
   ix35842 : inv02 port map ( Y=>nx35843, A=>nx34737);
   ix35844 : inv02 port map ( Y=>nx35845, A=>nx34737);
   ix35846 : inv02 port map ( Y=>nx35847, A=>nx34737);
   ix35848 : inv01 port map ( Y=>nx35849, A=>nx34821);
   ix35850 : inv02 port map ( Y=>nx35851, A=>nx35849);
   ix35852 : inv02 port map ( Y=>nx35853, A=>nx35849);
   ix35854 : inv02 port map ( Y=>nx35855, A=>nx35849);
   ix35856 : inv02 port map ( Y=>nx35857, A=>nx35849);
   ix35858 : inv02 port map ( Y=>nx35859, A=>nx35849);
   ix35860 : inv02 port map ( Y=>nx35861, A=>nx9490);
   ix35862 : inv02 port map ( Y=>nx35863, A=>nx9490);
   ix35864 : inv02 port map ( Y=>nx35865, A=>nx9490);
   ix35866 : inv01 port map ( Y=>nx35867, A=>nx34905);
   ix35868 : inv02 port map ( Y=>nx35869, A=>nx35867);
   ix35870 : inv02 port map ( Y=>nx35871, A=>nx35867);
   ix35872 : inv02 port map ( Y=>nx35873, A=>nx35867);
   ix35874 : inv01 port map ( Y=>nx35875, A=>nx34913);
   ix35876 : inv02 port map ( Y=>nx35877, A=>nx35875);
   ix35878 : inv02 port map ( Y=>nx35879, A=>nx35875);
   ix35880 : inv02 port map ( Y=>nx35881, A=>nx35875);
   ix35882 : inv02 port map ( Y=>nx35883, A=>nx35875);
   ix35884 : inv02 port map ( Y=>nx35885, A=>nx35875);
   ix35886 : inv02 port map ( Y=>nx35887, A=>nx12690);
   ix35888 : inv02 port map ( Y=>nx35889, A=>nx12690);
   ix35890 : inv02 port map ( Y=>nx35891, A=>nx12690);
   ix35892 : inv02 port map ( Y=>nx35893, A=>nx15874);
   ix35894 : inv02 port map ( Y=>nx35895, A=>nx15874);
   ix35896 : inv02 port map ( Y=>nx35897, A=>nx15874);
   ix35898 : inv02 port map ( Y=>nx35899, A=>nx17138);
   ix35900 : inv02 port map ( Y=>nx35901, A=>nx17138);
   ix35902 : inv02 port map ( Y=>nx35903, A=>nx17138);
   ix35904 : inv02 port map ( Y=>nx35905, A=>nx13373);
   ix35906 : inv02 port map ( Y=>nx35907, A=>nx13373);
   ix35908 : inv02 port map ( Y=>nx35909, A=>nx13373);
   ix35910 : inv02 port map ( Y=>nx35911, A=>done);
   ix35912 : inv02 port map ( Y=>nx35913, A=>done);
   ix35914 : inv02 port map ( Y=>nx35915, A=>done);
   ix35916 : inv02 port map ( Y=>nx35917, A=>done);
   ix35918 : inv02 port map ( Y=>nx35919, A=>nx36307);
   ix35920 : inv02 port map ( Y=>nx35921, A=>nx36307);
   ix35922 : inv02 port map ( Y=>nx35923, A=>nx36307);
   ix35924 : inv02 port map ( Y=>nx35925, A=>nx36309);
   ix35926 : inv02 port map ( Y=>nx35927, A=>nx36309);
   ix35928 : inv02 port map ( Y=>nx35929, A=>nx36309);
   ix35930 : inv02 port map ( Y=>nx35931, A=>nx36309);
   ix35932 : inv02 port map ( Y=>nx35933, A=>nx36309);
   ix35934 : inv02 port map ( Y=>nx35935, A=>nx36309);
   ix35936 : inv02 port map ( Y=>nx35937, A=>nx36309);
   ix35938 : inv02 port map ( Y=>nx35939, A=>nx36311);
   ix35940 : inv02 port map ( Y=>nx35941, A=>nx36311);
   ix35942 : inv02 port map ( Y=>nx35943, A=>nx36311);
   ix35944 : inv02 port map ( Y=>nx35945, A=>nx36311);
   ix35946 : inv02 port map ( Y=>nx35947, A=>nx36311);
   ix35948 : inv02 port map ( Y=>nx35949, A=>nx36311);
   ix35950 : inv02 port map ( Y=>nx35951, A=>nx36311);
   ix35952 : inv02 port map ( Y=>nx35953, A=>nx36313);
   ix35954 : inv02 port map ( Y=>nx35955, A=>nx36313);
   ix35956 : inv02 port map ( Y=>nx35957, A=>nx36313);
   ix35958 : inv02 port map ( Y=>nx35959, A=>nx36301);
   ix35960 : inv02 port map ( Y=>nx35961, A=>nx36301);
   ix35962 : inv02 port map ( Y=>nx35963, A=>nx36301);
   ix35964 : inv02 port map ( Y=>nx35965, A=>nx36301);
   ix35966 : inv02 port map ( Y=>nx35967, A=>nx36301);
   ix35968 : inv02 port map ( Y=>nx35969, A=>nx36301);
   ix35970 : inv02 port map ( Y=>nx35971, A=>nx36301);
   ix35972 : inv02 port map ( Y=>nx35973, A=>nx35735);
   ix35974 : inv02 port map ( Y=>nx35975, A=>nx35735);
   ix35976 : inv02 port map ( Y=>nx35977, A=>nx36331);
   ix35978 : inv02 port map ( Y=>nx35979, A=>nx36331);
   ix35980 : inv02 port map ( Y=>nx35981, A=>nx36331);
   ix35982 : inv02 port map ( Y=>nx35983, A=>nx36331);
   ix35984 : inv02 port map ( Y=>nx35985, A=>nx36333);
   ix35986 : inv02 port map ( Y=>nx35987, A=>nx36333);
   ix35988 : inv02 port map ( Y=>nx35989, A=>nx36333);
   ix35990 : inv02 port map ( Y=>nx35991, A=>nx36333);
   ix35992 : inv02 port map ( Y=>nx35993, A=>nx36333);
   ix35994 : inv02 port map ( Y=>nx35995, A=>nx36333);
   ix35996 : inv02 port map ( Y=>nx35997, A=>nx36333);
   ix35998 : inv02 port map ( Y=>nx35999, A=>nx36335);
   ix36000 : inv02 port map ( Y=>nx36001, A=>nx36335);
   ix36002 : inv02 port map ( Y=>nx36003, A=>nx36327);
   ix36004 : inv02 port map ( Y=>nx36005, A=>nx36327);
   ix36006 : inv02 port map ( Y=>nx36007, A=>nx36329);
   ix36008 : inv02 port map ( Y=>nx36009, A=>nx36329);
   ix36010 : inv02 port map ( Y=>nx36011, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix36012 : inv02 port map ( Y=>nx36013, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix36014 : inv02 port map ( Y=>nx36015, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix36016 : inv02 port map ( Y=>nx36017, A=>
      booth_booth_integrtaion_0_shift_reg_output_0);
   ix36018 : inv01 port map ( Y=>nx36019, A=>nx35289);
   ix36020 : inv02 port map ( Y=>nx36021, A=>nx36019);
   ix36022 : inv02 port map ( Y=>nx36023, A=>nx36019);
   ix36024 : inv02 port map ( Y=>nx36025, A=>nx36019);
   ix36026 : inv02 port map ( Y=>nx36027, A=>nx36019);
   ix36028 : inv02 port map ( Y=>nx36029, A=>nx36019);
   ix36030 : inv02 port map ( Y=>nx36031, A=>nx36341);
   ix36032 : inv02 port map ( Y=>nx36033, A=>nx36341);
   ix36034 : inv02 port map ( Y=>nx36035, A=>nx36343);
   ix36036 : inv02 port map ( Y=>nx36037, A=>nx36343);
   ix36038 : inv02 port map ( Y=>nx36039, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix36040 : inv02 port map ( Y=>nx36041, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix36042 : inv02 port map ( Y=>nx36043, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix36044 : inv02 port map ( Y=>nx36045, A=>
      booth_booth_integrtaion_8_shift_reg_output_0);
   ix36046 : inv02 port map ( Y=>nx36047, A=>nx36345);
   ix36048 : inv02 port map ( Y=>nx36049, A=>nx36345);
   ix36050 : inv02 port map ( Y=>nx36051, A=>nx36347);
   ix36052 : inv02 port map ( Y=>nx36053, A=>nx36347);
   ix36054 : inv02 port map ( Y=>nx36055, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix36056 : inv02 port map ( Y=>nx36057, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix36058 : inv02 port map ( Y=>nx36059, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix36060 : inv02 port map ( Y=>nx36061, A=>
      booth_booth_integrtaion_9_shift_reg_output_0);
   ix36062 : inv02 port map ( Y=>nx36063, A=>nx36337);
   ix36064 : inv02 port map ( Y=>nx36065, A=>nx36337);
   ix36066 : inv02 port map ( Y=>nx36067, A=>nx36339);
   ix36068 : inv02 port map ( Y=>nx36069, A=>nx36339);
   ix36070 : inv02 port map ( Y=>nx36071, A=>nx36339);
   ix36072 : inv02 port map ( Y=>nx36073, A=>nx36339);
   ix36074 : inv02 port map ( Y=>nx36075, A=>nx36339);
   ix36076 : inv02 port map ( Y=>nx36077, A=>nx36323);
   ix36078 : inv02 port map ( Y=>nx36079, A=>nx36323);
   ix36080 : inv02 port map ( Y=>nx36081, A=>nx36325);
   ix36082 : inv02 port map ( Y=>nx36083, A=>nx36325);
   ix36084 : inv02 port map ( Y=>nx36085, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix36086 : inv02 port map ( Y=>nx36087, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix36088 : inv02 port map ( Y=>nx36089, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix36090 : inv02 port map ( Y=>nx36091, A=>
      booth_booth_integrtaion_1_shift_reg_output_0);
   ix36092 : inv02 port map ( Y=>nx36093, A=>nx36319);
   ix36094 : inv02 port map ( Y=>nx36095, A=>nx36319);
   ix36096 : inv02 port map ( Y=>nx36097, A=>nx36321);
   ix36098 : inv02 port map ( Y=>nx36099, A=>nx36321);
   ix36100 : inv02 port map ( Y=>nx36101, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix36102 : inv02 port map ( Y=>nx36103, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix36104 : inv02 port map ( Y=>nx36105, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix36106 : inv02 port map ( Y=>nx36107, A=>
      booth_booth_integrtaion_2_shift_reg_output_0);
   ix36108 : inv02 port map ( Y=>nx36109, A=>nx36349);
   ix36110 : inv02 port map ( Y=>nx36111, A=>nx36349);
   ix36112 : inv02 port map ( Y=>nx36113, A=>nx36351);
   ix36114 : inv02 port map ( Y=>nx36115, A=>nx36351);
   ix36116 : inv02 port map ( Y=>nx36117, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix36118 : inv02 port map ( Y=>nx36119, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix36120 : inv02 port map ( Y=>nx36121, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix36122 : inv02 port map ( Y=>nx36123, A=>
      booth_booth_integrtaion_4_shift_reg_output_0);
   ix36124 : inv02 port map ( Y=>nx36125, A=>nx29498);
   ix36126 : inv02 port map ( Y=>nx36127, A=>nx29498);
   ix36128 : inv02 port map ( Y=>nx36129, A=>nx29498);
   ix36130 : inv02 port map ( Y=>nx36131, A=>nx36353);
   ix36132 : inv02 port map ( Y=>nx36133, A=>nx36353);
   ix36134 : inv02 port map ( Y=>nx36135, A=>nx36355);
   ix36136 : inv02 port map ( Y=>nx36137, A=>nx36355);
   ix36138 : inv02 port map ( Y=>nx36139, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix36140 : inv02 port map ( Y=>nx36141, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix36142 : inv02 port map ( Y=>nx36143, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix36144 : inv02 port map ( Y=>nx36145, A=>
      booth_booth_integrtaion_5_shift_reg_output_0);
   ix36146 : inv02 port map ( Y=>nx36147, A=>nx36315);
   ix36148 : inv02 port map ( Y=>nx36149, A=>nx36315);
   ix36150 : inv02 port map ( Y=>nx36151, A=>nx36317);
   ix36152 : inv02 port map ( Y=>nx36153, A=>nx36317);
   ix36154 : inv02 port map ( Y=>nx36155, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix36156 : inv02 port map ( Y=>nx36157, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix36158 : inv02 port map ( Y=>nx36159, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix36160 : inv02 port map ( Y=>nx36161, A=>
      booth_booth_integrtaion_3_shift_reg_output_0);
   ix36162 : inv02 port map ( Y=>nx36163, A=>nx36357);
   ix36164 : inv02 port map ( Y=>nx36165, A=>nx36357);
   ix36166 : inv02 port map ( Y=>nx36167, A=>nx36359);
   ix36168 : inv02 port map ( Y=>nx36169, A=>nx36359);
   ix36170 : inv02 port map ( Y=>nx36171, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix36172 : inv02 port map ( Y=>nx36173, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix36174 : inv02 port map ( Y=>nx36175, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix36176 : inv02 port map ( Y=>nx36177, A=>
      booth_booth_integrtaion_6_shift_reg_output_0);
   ix36178 : inv02 port map ( Y=>nx36179, A=>nx36361);
   ix36180 : inv02 port map ( Y=>nx36181, A=>nx36361);
   ix36182 : inv02 port map ( Y=>nx36183, A=>nx36363);
   ix36184 : inv02 port map ( Y=>nx36185, A=>nx36363);
   ix36186 : inv02 port map ( Y=>nx36187, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix36188 : inv02 port map ( Y=>nx36189, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix36190 : inv02 port map ( Y=>nx36191, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix36192 : inv02 port map ( Y=>nx36193, A=>
      booth_booth_integrtaion_7_shift_reg_output_0);
   ix36194 : inv02 port map ( Y=>nx36195, A=>nx29498);
   ix36196 : inv02 port map ( Y=>nx36197, A=>nx29498);
   ix36198 : inv02 port map ( Y=>nx36199, A=>nx29498);
   ix36200 : inv02 port map ( Y=>nx36201, A=>nx36365);
   ix36202 : inv02 port map ( Y=>nx36203, A=>nx36365);
   ix36204 : inv02 port map ( Y=>nx36205, A=>nx36365);
   ix36206 : inv02 port map ( Y=>nx36207, A=>nx36365);
   ix36208 : inv02 port map ( Y=>nx36209, A=>nx36367);
   ix36210 : inv02 port map ( Y=>nx36211, A=>nx36367);
   ix36212 : inv02 port map ( Y=>nx36213, A=>nx36367);
   ix36214 : inv02 port map ( Y=>nx36215, A=>nx36367);
   ix36216 : inv02 port map ( Y=>nx36217, A=>nx36367);
   ix36218 : inv02 port map ( Y=>nx36219, A=>nx36367);
   ix36220 : inv02 port map ( Y=>nx36221, A=>nx36367);
   ix36222 : inv02 port map ( Y=>nx36223, A=>nx36369);
   ix36224 : inv02 port map ( Y=>nx36225, A=>nx36369);
   ix36226 : inv02 port map ( Y=>nx36227, A=>nx36369);
   ix36228 : inv02 port map ( Y=>nx36229, A=>nx36369);
   ix36230 : inv02 port map ( Y=>nx36231, A=>nx36369);
   ix36232 : inv02 port map ( Y=>nx36233, A=>nx36369);
   ix36234 : inv02 port map ( Y=>nx36235, A=>nx36369);
   ix36236 : inv02 port map ( Y=>nx36237, A=>nx36371);
   ix36238 : inv02 port map ( Y=>nx36239, A=>nx36371);
   ix36240 : inv02 port map ( Y=>nx36241, A=>nx36373);
   ix36242 : inv02 port map ( Y=>nx36243, A=>nx36373);
   ix36244 : inv02 port map ( Y=>nx36245, A=>nx36373);
   ix36246 : inv02 port map ( Y=>nx36247, A=>nx36373);
   ix36248 : inv02 port map ( Y=>nx36249, A=>nx36375);
   ix36250 : inv02 port map ( Y=>nx36251, A=>nx36375);
   ix36252 : inv02 port map ( Y=>nx36253, A=>nx36375);
   ix36254 : inv02 port map ( Y=>nx36255, A=>nx36375);
   ix36256 : inv02 port map ( Y=>nx36257, A=>nx36375);
   ix36258 : inv02 port map ( Y=>nx36259, A=>nx36375);
   ix36260 : inv02 port map ( Y=>nx36261, A=>nx36375);
   ix36262 : inv02 port map ( Y=>nx36263, A=>nx36377);
   ix36264 : inv02 port map ( Y=>nx36265, A=>nx36377);
   ix36266 : inv02 port map ( Y=>nx36267, A=>nx36377);
   ix36268 : inv02 port map ( Y=>nx36269, A=>nx36377);
   ix36270 : inv02 port map ( Y=>nx36271, A=>nx36377);
   ix36272 : inv02 port map ( Y=>nx36273, A=>nx36377);
   ix36274 : inv02 port map ( Y=>nx36275, A=>nx36377);
   ix36276 : inv02 port map ( Y=>nx36277, A=>nx36379);
   ix36278 : inv02 port map ( Y=>nx36279, A=>nx36379);
   ix36280 : inv02 port map ( Y=>nx36281, A=>nx36385);
   ix36282 : inv02 port map ( Y=>nx36283, A=>nx36385);
   ix36284 : inv02 port map ( Y=>nx36285, A=>nx36385);
   ix36286 : inv02 port map ( Y=>nx36287, A=>nx36385);
   ix36288 : inv02 port map ( Y=>nx36289, A=>nx36385);
   ix36290 : inv02 port map ( Y=>nx36291, A=>nx36381);
   ix36292 : inv02 port map ( Y=>nx36293, A=>nx36381);
   ix36294 : inv02 port map ( Y=>nx36295, A=>nx36381);
   ix36296 : inv02 port map ( Y=>nx36297, A=>nx36383);
   ix36298 : inv02 port map ( Y=>nx36299, A=>nx35173);
   ix36300 : inv02 port map ( Y=>nx36301, A=>nx35173);
   ix36306 : inv02 port map ( Y=>nx36307, A=>nx35163);
   ix36308 : inv02 port map ( Y=>nx36309, A=>nx35163);
   ix36310 : inv02 port map ( Y=>nx36311, A=>nx35163);
   ix36312 : inv02 port map ( Y=>nx36313, A=>nx35163);
   ix36314 : inv02 port map ( Y=>nx36315, A=>nx35499);
   ix36316 : inv02 port map ( Y=>nx36317, A=>nx35499);
   ix36318 : inv02 port map ( Y=>nx36319, A=>nx35399);
   ix36320 : inv02 port map ( Y=>nx36321, A=>nx35399);
   ix36322 : inv02 port map ( Y=>nx36323, A=>nx35373);
   ix36324 : inv02 port map ( Y=>nx36325, A=>nx35373);
   ix36326 : inv02 port map ( Y=>nx36327, A=>nx35193);
   ix36328 : inv02 port map ( Y=>nx36329, A=>nx35193);
   ix36330 : inv02 port map ( Y=>nx36331, A=>nx35187);
   ix36332 : inv02 port map ( Y=>nx36333, A=>nx35187);
   ix36334 : inv02 port map ( Y=>nx36335, A=>nx35187);
   ix36336 : inv02 port map ( Y=>nx36337, A=>nx36385);
   ix36338 : inv02 port map ( Y=>nx36339, A=>nx36385);
   ix36340 : inv02 port map ( Y=>nx36341, A=>nx35301);
   ix36342 : inv02 port map ( Y=>nx36343, A=>nx35301);
   ix36344 : inv02 port map ( Y=>nx36345, A=>nx35327);
   ix36346 : inv02 port map ( Y=>nx36347, A=>nx35327);
   ix36348 : inv02 port map ( Y=>nx36349, A=>nx35425);
   ix36350 : inv02 port map ( Y=>nx36351, A=>nx35425);
   ix36352 : inv02 port map ( Y=>nx36353, A=>nx35473);
   ix36354 : inv02 port map ( Y=>nx36355, A=>nx35473);
   ix36356 : inv02 port map ( Y=>nx36357, A=>nx35525);
   ix36358 : inv02 port map ( Y=>nx36359, A=>nx35525);
   ix36360 : inv02 port map ( Y=>nx36361, A=>nx35551);
   ix36362 : inv02 port map ( Y=>nx36363, A=>nx35551);
   ix36364 : inv02 port map ( Y=>nx36365, A=>nx35595);
   ix36366 : inv02 port map ( Y=>nx36367, A=>nx35595);
   ix36368 : inv02 port map ( Y=>nx36369, A=>nx35595);
   ix36370 : inv02 port map ( Y=>nx36371, A=>nx35595);
   ix36372 : inv02 port map ( Y=>nx36373, A=>nx35603);
   ix36374 : inv02 port map ( Y=>nx36375, A=>nx35603);
   ix36376 : inv02 port map ( Y=>nx36377, A=>nx35603);
   ix36378 : inv02 port map ( Y=>nx36379, A=>nx35603);
   ix36380 : inv02 port map ( Y=>nx36381, A=>nx35747);
   ix36382 : inv02 port map ( Y=>nx36383, A=>nx35747);
   ix36384 : inv02 port map ( Y=>nx36385, A=>nx6352);
   ix36386 : inv02 port map ( Y=>nx36387, A=>enable_decoder_dst_booth);
   ix36388 : inv02 port map ( Y=>nx36389, A=>max_calc_state_2);
   ix36390 : inv02 port map ( Y=>nx36391, A=>nx26669);
   ix36392 : inv02 port map ( Y=>nx36393, A=>nx26675);
end a_controller ;

