
-- 
-- Definition of  booth_adder_components
-- 
--      Fri Apr 19 17:55:29 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.adk_components.all;

entity booth_adder_components is
   port (
      clk : IN std_logic ;
      rst : IN std_logic ;
      set : IN std_logic ;
      done : OUT std_logic ;
      neuron : IN std_logic_vector (15 DOWNTO 0) ;
      weight_0 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_1 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_2 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_3 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_4 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_5 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_6 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_7 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_8 : IN std_logic_vector (15 DOWNTO 0) ;
      weight_9 : IN std_logic_vector (15 DOWNTO 0) ;
      label_0 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_1 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_2 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_3 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_4 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_5 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_6 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_7 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_8 : OUT std_logic_vector (15 DOWNTO 0) ;
      label_9 : OUT std_logic_vector (15 DOWNTO 0) ;
      adderInput_0 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_1 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_2 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_3 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_4 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_5 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_6 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_7 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_8 : IN std_logic_vector (15 DOWNTO 0) ;
      adderInput_9 : IN std_logic_vector (15 DOWNTO 0) ;
      dec_enable : OUT std_logic ;
      dec_sel : OUT std_logic_vector (3 DOWNTO 0)) ;
end booth_adder_components ;

architecture my_booth_adder_components of booth_adder_components is
   signal dec_sel_0_EXMPLR, booth_integration_output_9_0, 
      booth_integrtaion_9_shift_reg_output_9, 
      booth_integrtaion_9_shift_Reg_count_9, 
      booth_integrtaion_9_shift_Reg_output_8, 
      booth_integrtaion_9_shift_Reg_count_8, 
      booth_integrtaion_9_shift_Reg_output_7, 
      booth_integrtaion_9_shift_Reg_count_7, 
      booth_integrtaion_9_shift_Reg_output_6, 
      booth_integrtaion_9_shift_Reg_count_6, 
      booth_integrtaion_9_shift_Reg_output_5, 
      booth_integrtaion_9_shift_Reg_count_5, 
      booth_integrtaion_9_shift_Reg_output_4, 
      booth_integrtaion_9_shift_Reg_count_4, 
      booth_integrtaion_9_shift_Reg_output_3, 
      booth_integrtaion_9_shift_Reg_count_3, 
      booth_integrtaion_9_shift_Reg_output_2, 
      booth_integrtaion_9_shift_Reg_count_2, 
      booth_integrtaion_9_shift_Reg_output_1, 
      booth_integrtaion_9_shift_Reg_count_1, 
      booth_integrtaion_9_shift_reg_output_0, 
      booth_integrtaion_9_shift_Reg_count_0, booth_integration_output_9_1, 
      booth_integration_output_9_2, booth_integration_output_9_3, 
      booth_integration_output_9_4, booth_integration_output_9_5, 
      booth_integration_output_9_6, booth_integration_output_9_7, 
      booth_integration_output_9_8, booth_integration_output_9_9, 
      booth_integration_output_9_10, booth_integration_output_9_11, 
      booth_integration_output_9_12, booth_integration_output_9_13, 
      booth_integration_output_9_14, booth_integration_output_9_15, 
      booth_integrtaion_9_booth_output_16, nx102, nx106, nx112, 
      booth_integrtaion_9_booth_output_17, nx2805, nx120, nx136, nx2807, 
      nx146, nx150, nx164, booth_integrtaion_9_booth_output_19, nx2808, 
      nx174, nx184, nx198, nx208, nx212, booth_integrtaion_9_booth_output_21, 
      nx2810, nx222, nx232, nx246, nx256, nx260, 
      booth_integrtaion_9_booth_output_23, nx2813, nx270, nx280, nx294, 
      nx304, nx308, booth_integrtaion_9_booth_output_25, nx2817, nx318, 
      nx328, nx342, nx352, nx356, booth_integrtaion_9_booth_output_27, 
      nx2821, nx366, nx376, nx390, nx400, nx404, 
      booth_integrtaion_9_booth_output_29, nx2825, nx414, nx424, 
      booth_integrtaion_9_booth_output_31, nx438, nx448, nx452, nx454, nx462, 
      nx468, nx480, nx488, nx504, nx512, nx528, nx536, nx552, nx560, nx576, 
      nx584, nx600, nx608, nx620, nx636, nx642, nx648, nx666, nx678, nx690, 
      nx702, nx714, nx726, nx738, nx750, nx762, nx774, nx786, nx798, nx810, 
      nx822, nx834, nx842, nx856, nx858, nx872, nx874, nx888, nx890, nx904, 
      nx906, nx920, nx922, nx936, nx938, nx952, booth_integration_output_8_0, 
      booth_integrtaion_8_shift_reg_output_9, 
      booth_integrtaion_8_shift_Reg_count_9, 
      booth_integrtaion_8_shift_Reg_output_8, 
      booth_integrtaion_8_shift_Reg_count_8, 
      booth_integrtaion_8_shift_Reg_output_7, 
      booth_integrtaion_8_shift_Reg_count_7, 
      booth_integrtaion_8_shift_Reg_output_6, 
      booth_integrtaion_8_shift_Reg_count_6, 
      booth_integrtaion_8_shift_Reg_output_5, 
      booth_integrtaion_8_shift_Reg_count_5, 
      booth_integrtaion_8_shift_Reg_output_4, 
      booth_integrtaion_8_shift_Reg_count_4, 
      booth_integrtaion_8_shift_Reg_output_3, 
      booth_integrtaion_8_shift_Reg_count_3, 
      booth_integrtaion_8_shift_Reg_output_2, 
      booth_integrtaion_8_shift_Reg_count_2, 
      booth_integrtaion_8_shift_Reg_output_1, 
      booth_integrtaion_8_shift_Reg_count_1, 
      booth_integrtaion_8_shift_reg_output_0, 
      booth_integrtaion_8_shift_Reg_count_0, booth_integration_output_8_1, 
      booth_integration_output_8_2, booth_integration_output_8_3, 
      booth_integration_output_8_4, booth_integration_output_8_5, 
      booth_integration_output_8_6, booth_integration_output_8_7, 
      booth_integration_output_8_8, booth_integration_output_8_9, 
      booth_integration_output_8_10, booth_integration_output_8_11, 
      booth_integration_output_8_12, booth_integration_output_8_13, 
      booth_integration_output_8_14, booth_integration_output_8_15, 
      booth_integrtaion_8_booth_output_16, nx1088, nx1092, nx1098, 
      booth_integrtaion_8_booth_output_17, nx2831, nx1106, nx1122, nx2833, 
      nx1132, nx1136, nx1150, booth_integrtaion_8_booth_output_19, nx2835, 
      nx1160, nx1170, nx1184, nx1194, nx1198, 
      booth_integrtaion_8_booth_output_21, nx2839, nx1208, nx1218, nx1232, 
      nx1242, nx1246, booth_integrtaion_8_booth_output_23, nx2843, nx1256, 
      nx1266, nx1280, nx1290, nx1294, booth_integrtaion_8_booth_output_25, 
      nx2847, nx1304, nx1314, nx1328, nx1338, nx1342, 
      booth_integrtaion_8_booth_output_27, nx2851, nx1352, nx1362, nx1376, 
      nx1386, nx1390, booth_integrtaion_8_booth_output_29, nx2855, nx1400, 
      nx1410, booth_integrtaion_8_booth_output_31, nx1424, nx1434, nx1438, 
      nx1440, nx1448, nx1454, nx1466, nx1474, nx1490, nx1498, nx1514, nx1522, 
      nx1538, nx1546, nx1562, nx1570, nx1586, nx1594, nx1606, nx1622, nx1628, 
      nx1634, nx1652, nx1664, nx1676, nx1688, nx1700, nx1712, nx1724, nx1736, 
      nx1748, nx1760, nx1772, nx1784, nx1796, nx1808, nx1820, nx1828, nx1842, 
      nx1844, nx1858, nx1860, nx1874, nx1876, nx1890, nx1892, nx1906, nx1908, 
      nx1922, nx1924, nx1938, booth_integration_output_7_0, 
      booth_integrtaion_7_shift_reg_output_9, 
      booth_integrtaion_7_shift_Reg_count_9, 
      booth_integrtaion_7_shift_Reg_output_8, 
      booth_integrtaion_7_shift_Reg_count_8, 
      booth_integrtaion_7_shift_Reg_output_7, 
      booth_integrtaion_7_shift_Reg_count_7, 
      booth_integrtaion_7_shift_Reg_output_6, 
      booth_integrtaion_7_shift_Reg_count_6, 
      booth_integrtaion_7_shift_Reg_output_5, 
      booth_integrtaion_7_shift_Reg_count_5, 
      booth_integrtaion_7_shift_Reg_output_4, 
      booth_integrtaion_7_shift_Reg_count_4, 
      booth_integrtaion_7_shift_Reg_output_3, 
      booth_integrtaion_7_shift_Reg_count_3, 
      booth_integrtaion_7_shift_Reg_output_2, 
      booth_integrtaion_7_shift_Reg_count_2, 
      booth_integrtaion_7_shift_Reg_output_1, 
      booth_integrtaion_7_shift_Reg_count_1, 
      booth_integrtaion_7_shift_reg_output_0, 
      booth_integrtaion_7_shift_Reg_count_0, booth_integration_output_7_1, 
      booth_integration_output_7_2, booth_integration_output_7_3, 
      booth_integration_output_7_4, booth_integration_output_7_5, 
      booth_integration_output_7_6, booth_integration_output_7_7, 
      booth_integration_output_7_8, booth_integration_output_7_9, 
      booth_integration_output_7_10, booth_integration_output_7_11, 
      booth_integration_output_7_12, booth_integration_output_7_13, 
      booth_integration_output_7_14, booth_integration_output_7_15, 
      booth_integrtaion_7_booth_output_16, nx2074, nx2078, nx2084, 
      booth_integrtaion_7_booth_output_17, nx2861, nx2092, nx2108, nx2863, 
      nx2118, nx2122, nx2136, booth_integrtaion_7_booth_output_19, nx2865, 
      nx2146, nx2156, nx2170, nx2180, nx2184, 
      booth_integrtaion_7_booth_output_21, nx2869, nx2194, nx2204, nx2218, 
      nx2228, nx2232, booth_integrtaion_7_booth_output_23, nx2873, nx2242, 
      nx2252, nx2266, nx2276, nx2280, booth_integrtaion_7_booth_output_25, 
      nx2877, nx2290, nx2300, nx2314, nx2324, nx2328, 
      booth_integrtaion_7_booth_output_27, nx2881, nx2338, nx2348, nx2362, 
      nx2372, nx2376, booth_integrtaion_7_booth_output_29, nx2885, nx2386, 
      nx2396, booth_integrtaion_7_booth_output_31, nx2410, nx2420, nx2424, 
      nx2426, nx2434, nx2440, nx2452, nx2460, nx2476, nx2484, nx2500, nx2508, 
      nx2524, nx2532, nx2548, nx2556, nx2572, nx2580, nx2592, nx2608, nx2614, 
      nx2620, nx2638, nx2650, nx2662, nx2674, nx2686, nx2698, nx2710, nx2722, 
      nx2734, nx2746, nx2758, nx2770, nx2782, nx2794, nx2806, nx2814, nx2828, 
      nx2830, nx2844, nx2846, nx2860, nx2862, nx2876, nx2878, nx2892, nx2894, 
      nx2908, nx2910, nx2924, booth_integration_output_6_0, 
      booth_integrtaion_6_shift_reg_output_9, 
      booth_integrtaion_6_shift_Reg_count_9, 
      booth_integrtaion_6_shift_Reg_output_8, 
      booth_integrtaion_6_shift_Reg_count_8, 
      booth_integrtaion_6_shift_Reg_output_7, 
      booth_integrtaion_6_shift_Reg_count_7, 
      booth_integrtaion_6_shift_Reg_output_6, 
      booth_integrtaion_6_shift_Reg_count_6, 
      booth_integrtaion_6_shift_Reg_output_5, 
      booth_integrtaion_6_shift_Reg_count_5, 
      booth_integrtaion_6_shift_Reg_output_4, 
      booth_integrtaion_6_shift_Reg_count_4, 
      booth_integrtaion_6_shift_Reg_output_3, 
      booth_integrtaion_6_shift_Reg_count_3, 
      booth_integrtaion_6_shift_Reg_output_2, 
      booth_integrtaion_6_shift_Reg_count_2, 
      booth_integrtaion_6_shift_Reg_output_1, 
      booth_integrtaion_6_shift_Reg_count_1, 
      booth_integrtaion_6_shift_reg_output_0, 
      booth_integrtaion_6_shift_Reg_count_0, booth_integration_output_6_1, 
      booth_integration_output_6_2, booth_integration_output_6_3, 
      booth_integration_output_6_4, booth_integration_output_6_5, 
      booth_integration_output_6_6, booth_integration_output_6_7, 
      booth_integration_output_6_8, booth_integration_output_6_9, 
      booth_integration_output_6_10, booth_integration_output_6_11, 
      booth_integration_output_6_12, booth_integration_output_6_13, 
      booth_integration_output_6_14, booth_integration_output_6_15, 
      booth_integrtaion_6_booth_output_16, nx3060, nx3064, nx3070, 
      booth_integrtaion_6_booth_output_17, nx2891, nx3078, nx3094, nx2893, 
      nx3104, nx3108, nx3122, booth_integrtaion_6_booth_output_19, nx2895, 
      nx3132, nx3142, nx3156, nx3166, nx3170, 
      booth_integrtaion_6_booth_output_21, nx2899, nx3180, nx3190, nx3204, 
      nx3214, nx3218, booth_integrtaion_6_booth_output_23, nx2903, nx3228, 
      nx3238, nx3252, nx3262, nx3266, booth_integrtaion_6_booth_output_25, 
      nx2907, nx3276, nx3286, nx3300, nx3310, nx3314, 
      booth_integrtaion_6_booth_output_27, nx2911, nx3324, nx3334, nx3348, 
      nx3358, nx3362, booth_integrtaion_6_booth_output_29, nx2915, nx3372, 
      nx3382, booth_integrtaion_6_booth_output_31, nx3396, nx3406, nx3410, 
      nx3412, nx3420, nx3426, nx3438, nx3446, nx3462, nx3470, nx3486, nx3494, 
      nx3510, nx3518, nx3534, nx3542, nx3558, nx3566, nx3578, nx3594, nx3600, 
      nx3606, nx3624, nx3636, nx3648, nx3660, nx3672, nx3684, nx3696, nx3708, 
      nx3720, nx3732, nx3744, nx3756, nx3768, nx3780, nx3792, nx3800, nx3814, 
      nx3816, nx3830, nx3832, nx3846, nx3848, nx3862, nx3864, nx3878, nx3880, 
      nx3894, nx3896, nx3910, booth_integration_output_5_0, 
      booth_integrtaion_5_shift_reg_output_9, 
      booth_integrtaion_5_shift_Reg_count_9, 
      booth_integrtaion_5_shift_Reg_output_8, 
      booth_integrtaion_5_shift_Reg_count_8, 
      booth_integrtaion_5_shift_Reg_output_7, 
      booth_integrtaion_5_shift_Reg_count_7, 
      booth_integrtaion_5_shift_Reg_output_6, 
      booth_integrtaion_5_shift_Reg_count_6, 
      booth_integrtaion_5_shift_Reg_output_5, 
      booth_integrtaion_5_shift_Reg_count_5, 
      booth_integrtaion_5_shift_Reg_output_4, 
      booth_integrtaion_5_shift_Reg_count_4, 
      booth_integrtaion_5_shift_Reg_output_3, 
      booth_integrtaion_5_shift_Reg_count_3, 
      booth_integrtaion_5_shift_Reg_output_2, 
      booth_integrtaion_5_shift_Reg_count_2, 
      booth_integrtaion_5_shift_Reg_output_1, 
      booth_integrtaion_5_shift_Reg_count_1, 
      booth_integrtaion_5_shift_reg_output_0, 
      booth_integrtaion_5_shift_Reg_count_0, booth_integration_output_5_1, 
      booth_integration_output_5_2, booth_integration_output_5_3, 
      booth_integration_output_5_4, booth_integration_output_5_5, 
      booth_integration_output_5_6, booth_integration_output_5_7, 
      booth_integration_output_5_8, booth_integration_output_5_9, 
      booth_integration_output_5_10, booth_integration_output_5_11, 
      booth_integration_output_5_12, booth_integration_output_5_13, 
      booth_integration_output_5_14, booth_integration_output_5_15, 
      booth_integrtaion_5_booth_output_16, nx4046, nx4050, nx4056, 
      booth_integrtaion_5_booth_output_17, nx2921, nx4064, nx4080, nx2923, 
      nx4090, nx4094, nx4108, booth_integrtaion_5_booth_output_19, nx2925, 
      nx4118, nx4128, nx4142, nx4152, nx4156, 
      booth_integrtaion_5_booth_output_21, nx2928, nx4166, nx4176, nx4190, 
      nx4200, nx4204, booth_integrtaion_5_booth_output_23, nx2930, nx4214, 
      nx4224, nx4238, nx4248, nx4252, booth_integrtaion_5_booth_output_25, 
      nx2932, nx4262, nx4272, nx4286, nx4296, nx4300, 
      booth_integrtaion_5_booth_output_27, nx2934, nx4310, nx4320, nx4334, 
      nx4344, nx4348, booth_integrtaion_5_booth_output_29, nx2936, nx4358, 
      nx4368, booth_integrtaion_5_booth_output_31, nx4382, nx4392, nx4396, 
      nx4398, nx4406, nx4412, nx4424, nx4432, nx4448, nx4456, nx4472, nx4480, 
      nx4496, nx4504, nx4520, nx4528, nx4544, nx4552, nx4564, nx4580, nx4586, 
      nx4592, nx4610, nx4622, nx4634, nx4646, nx4658, nx4670, nx4682, nx4694, 
      nx4706, nx4718, nx4730, nx4742, nx4754, nx4766, nx4778, nx4786, nx4800, 
      nx4802, nx4816, nx4818, nx4832, nx4834, nx4848, nx4850, nx4864, nx4866, 
      nx4880, nx4882, nx4896, booth_integration_output_4_0, 
      booth_integrtaion_4_shift_reg_output_9, 
      booth_integrtaion_4_shift_Reg_count_9, 
      booth_integrtaion_4_shift_Reg_output_8, 
      booth_integrtaion_4_shift_Reg_count_8, 
      booth_integrtaion_4_shift_Reg_output_7, 
      booth_integrtaion_4_shift_Reg_count_7, 
      booth_integrtaion_4_shift_Reg_output_6, 
      booth_integrtaion_4_shift_Reg_count_6, 
      booth_integrtaion_4_shift_Reg_output_5, 
      booth_integrtaion_4_shift_Reg_count_5, 
      booth_integrtaion_4_shift_Reg_output_4, 
      booth_integrtaion_4_shift_Reg_count_4, 
      booth_integrtaion_4_shift_Reg_output_3, 
      booth_integrtaion_4_shift_Reg_count_3, 
      booth_integrtaion_4_shift_Reg_output_2, 
      booth_integrtaion_4_shift_Reg_count_2, 
      booth_integrtaion_4_shift_Reg_output_1, 
      booth_integrtaion_4_shift_Reg_count_1, 
      booth_integrtaion_4_shift_reg_output_0, 
      booth_integrtaion_4_shift_Reg_count_0, booth_integration_output_4_1, 
      booth_integration_output_4_2, booth_integration_output_4_3, 
      booth_integration_output_4_4, booth_integration_output_4_5, 
      booth_integration_output_4_6, booth_integration_output_4_7, 
      booth_integration_output_4_8, booth_integration_output_4_9, 
      booth_integration_output_4_10, booth_integration_output_4_11, 
      booth_integration_output_4_12, booth_integration_output_4_13, 
      booth_integration_output_4_14, booth_integration_output_4_15, 
      booth_integrtaion_4_booth_output_16, nx5032, nx5036, nx5042, 
      booth_integrtaion_4_booth_output_17, nx2939, nx5050, nx5066, nx2940, 
      nx5076, nx5080, nx5094, booth_integrtaion_4_booth_output_19, nx2941, 
      nx5104, nx5114, nx5128, nx5138, nx5142, 
      booth_integrtaion_4_booth_output_21, nx2943, nx5152, nx5162, nx5176, 
      nx5186, nx5190, booth_integrtaion_4_booth_output_23, nx2945, nx5200, 
      nx5210, nx5224, nx5234, nx5238, booth_integrtaion_4_booth_output_25, 
      nx2947, nx5248, nx5258, nx5272, nx5282, nx5286, 
      booth_integrtaion_4_booth_output_27, nx2949, nx5296, nx5306, nx5320, 
      nx5330, nx5334, booth_integrtaion_4_booth_output_29, nx2951, nx5344, 
      nx5354, booth_integrtaion_4_booth_output_31, nx5368, nx5378, nx5382, 
      nx5384, nx5392, nx5398, nx5410, nx5418, nx5434, nx5442, nx5458, nx5466, 
      nx5482, nx5490, nx5506, nx5514, nx5530, nx5538, nx5550, nx5566, nx5572, 
      nx5578, nx5596, nx5608, nx5620, nx5632, nx5644, nx5656, nx5668, nx5680, 
      nx5692, nx5704, nx5716, nx5728, nx5740, nx5752, nx5764, nx5772, nx5786, 
      nx5788, nx5802, nx5804, nx5818, nx5820, nx5834, nx5836, nx5850, nx5852, 
      nx5866, nx5868, nx5882, booth_integration_output_3_0, 
      booth_integrtaion_3_shift_reg_output_9, 
      booth_integrtaion_3_shift_Reg_count_9, 
      booth_integrtaion_3_shift_Reg_output_8, 
      booth_integrtaion_3_shift_Reg_count_8, 
      booth_integrtaion_3_shift_Reg_output_7, 
      booth_integrtaion_3_shift_Reg_count_7, 
      booth_integrtaion_3_shift_Reg_output_6, 
      booth_integrtaion_3_shift_Reg_count_6, 
      booth_integrtaion_3_shift_Reg_output_5, 
      booth_integrtaion_3_shift_Reg_count_5, 
      booth_integrtaion_3_shift_Reg_output_4, 
      booth_integrtaion_3_shift_Reg_count_4, 
      booth_integrtaion_3_shift_Reg_output_3, 
      booth_integrtaion_3_shift_Reg_count_3, 
      booth_integrtaion_3_shift_Reg_output_2, 
      booth_integrtaion_3_shift_Reg_count_2, 
      booth_integrtaion_3_shift_Reg_output_1, 
      booth_integrtaion_3_shift_Reg_count_1, 
      booth_integrtaion_3_shift_reg_output_0, 
      booth_integrtaion_3_shift_Reg_count_0, booth_integration_output_3_1, 
      booth_integration_output_3_2, booth_integration_output_3_3, 
      booth_integration_output_3_4, booth_integration_output_3_5, 
      booth_integration_output_3_6, booth_integration_output_3_7, 
      booth_integration_output_3_8, booth_integration_output_3_9, 
      booth_integration_output_3_10, booth_integration_output_3_11, 
      booth_integration_output_3_12, booth_integration_output_3_13, 
      booth_integration_output_3_14, booth_integration_output_3_15, 
      booth_integrtaion_3_booth_output_16, nx6018, nx6022, nx6028, 
      booth_integrtaion_3_booth_output_17, nx2954, nx6036, nx6052, nx2955, 
      nx6062, nx6066, nx6080, booth_integrtaion_3_booth_output_19, nx2956, 
      nx6090, nx6100, nx6114, nx6124, nx6128, 
      booth_integrtaion_3_booth_output_21, nx2959, nx6138, nx6148, nx6162, 
      nx6172, nx6176, booth_integrtaion_3_booth_output_23, nx2961, nx6186, 
      nx6196, nx6210, nx6220, nx6224, booth_integrtaion_3_booth_output_25, 
      nx2963, nx6234, nx6244, nx6258, nx6268, nx6272, 
      booth_integrtaion_3_booth_output_27, nx2965, nx6282, nx6292, nx6306, 
      nx6316, nx6320, booth_integrtaion_3_booth_output_29, nx2967, nx6330, 
      nx6340, booth_integrtaion_3_booth_output_31, nx6354, nx6364, nx6368, 
      nx6370, nx6378, nx6384, nx6396, nx6404, nx6420, nx6428, nx6444, nx6452, 
      nx6468, nx6476, nx6492, nx6500, nx6516, nx6524, nx6536, nx6552, nx6558, 
      nx6564, nx6582, nx6594, nx6606, nx6618, nx6630, nx6642, nx6654, nx6666, 
      nx6678, nx6690, nx6702, nx6714, nx6726, nx6738, nx6750, nx6758, nx6772, 
      nx6774, nx6788, nx6790, nx6804, nx6806, nx6820, nx6822, nx6836, nx6838, 
      nx6852, nx6854, nx6868, booth_integration_output_2_0, 
      booth_integrtaion_2_shift_reg_output_9, 
      booth_integrtaion_2_shift_Reg_count_9, 
      booth_integrtaion_2_shift_Reg_output_8, 
      booth_integrtaion_2_shift_Reg_count_8, 
      booth_integrtaion_2_shift_Reg_output_7, 
      booth_integrtaion_2_shift_Reg_count_7, 
      booth_integrtaion_2_shift_Reg_output_6, 
      booth_integrtaion_2_shift_Reg_count_6, 
      booth_integrtaion_2_shift_Reg_output_5, 
      booth_integrtaion_2_shift_Reg_count_5, 
      booth_integrtaion_2_shift_Reg_output_4, 
      booth_integrtaion_2_shift_Reg_count_4, 
      booth_integrtaion_2_shift_Reg_output_3, 
      booth_integrtaion_2_shift_Reg_count_3, 
      booth_integrtaion_2_shift_Reg_output_2, 
      booth_integrtaion_2_shift_Reg_count_2, 
      booth_integrtaion_2_shift_Reg_output_1, 
      booth_integrtaion_2_shift_Reg_count_1, 
      booth_integrtaion_2_shift_reg_output_0, 
      booth_integrtaion_2_shift_Reg_count_0, booth_integration_output_2_1, 
      booth_integration_output_2_2, booth_integration_output_2_3, 
      booth_integration_output_2_4, booth_integration_output_2_5, 
      booth_integration_output_2_6, booth_integration_output_2_7, 
      booth_integration_output_2_8, booth_integration_output_2_9, 
      booth_integration_output_2_10, booth_integration_output_2_11, 
      booth_integration_output_2_12, booth_integration_output_2_13, 
      booth_integration_output_2_14, booth_integration_output_2_15, 
      booth_integrtaion_2_booth_output_16, nx7004, nx7008, nx7014, 
      booth_integrtaion_2_booth_output_17, nx2970, nx7022, nx7038, nx2971, 
      nx7048, nx7052, nx7066, booth_integrtaion_2_booth_output_19, nx2972, 
      nx7076, nx7086, nx7100, nx7110, nx7114, 
      booth_integrtaion_2_booth_output_21, nx2974, nx7124, nx7134, nx7148, 
      nx7158, nx7162, booth_integrtaion_2_booth_output_23, nx2976, nx7172, 
      nx7182, nx7196, nx7206, nx7210, booth_integrtaion_2_booth_output_25, 
      nx2978, nx7220, nx7230, nx7244, nx7254, nx7258, 
      booth_integrtaion_2_booth_output_27, nx2980, nx7268, nx7278, nx7292, 
      nx7302, nx7306, booth_integrtaion_2_booth_output_29, nx2982, nx7316, 
      nx7326, booth_integrtaion_2_booth_output_31, nx7340, nx7350, nx7354, 
      nx7356, nx7364, nx7370, nx7382, nx7390, nx7406, nx7414, nx7430, nx7438, 
      nx7454, nx7462, nx7478, nx7486, nx7502, nx7510, nx7522, nx7538, nx7544, 
      nx7550, nx7568, nx7580, nx7592, nx7604, nx7616, nx7628, nx7640, nx7652, 
      nx7664, nx7676, nx7688, nx7700, nx7712, nx7724, nx7736, nx7744, nx7758, 
      nx7760, nx7774, nx7776, nx7790, nx7792, nx7806, nx7808, nx7822, nx7824, 
      nx7838, nx7840, nx7854, booth_integration_output_1_0, 
      booth_integrtaion_1_shift_reg_output_9, 
      booth_integrtaion_1_shift_Reg_count_9, 
      booth_integrtaion_1_shift_Reg_output_8, 
      booth_integrtaion_1_shift_Reg_count_8, 
      booth_integrtaion_1_shift_Reg_output_7, 
      booth_integrtaion_1_shift_Reg_count_7, 
      booth_integrtaion_1_shift_Reg_output_6, 
      booth_integrtaion_1_shift_Reg_count_6, 
      booth_integrtaion_1_shift_Reg_output_5, 
      booth_integrtaion_1_shift_Reg_count_5, 
      booth_integrtaion_1_shift_Reg_output_4, 
      booth_integrtaion_1_shift_Reg_count_4, 
      booth_integrtaion_1_shift_Reg_output_3, 
      booth_integrtaion_1_shift_Reg_count_3, 
      booth_integrtaion_1_shift_Reg_output_2, 
      booth_integrtaion_1_shift_Reg_count_2, 
      booth_integrtaion_1_shift_Reg_output_1, 
      booth_integrtaion_1_shift_Reg_count_1, 
      booth_integrtaion_1_shift_reg_output_0, 
      booth_integrtaion_1_shift_Reg_count_0, booth_integration_output_1_1, 
      booth_integration_output_1_2, booth_integration_output_1_3, 
      booth_integration_output_1_4, booth_integration_output_1_5, 
      booth_integration_output_1_6, booth_integration_output_1_7, 
      booth_integration_output_1_8, booth_integration_output_1_9, 
      booth_integration_output_1_10, booth_integration_output_1_11, 
      booth_integration_output_1_12, booth_integration_output_1_13, 
      booth_integration_output_1_14, booth_integration_output_1_15, 
      booth_integrtaion_1_booth_output_16, nx7990, nx7994, nx8000, 
      booth_integrtaion_1_booth_output_17, nx2985, nx8008, nx8024, nx2986, 
      nx8034, nx8038, nx8052, booth_integrtaion_1_booth_output_19, nx2987, 
      nx8062, nx8072, nx8086, nx8096, nx8100, 
      booth_integrtaion_1_booth_output_21, nx2989, nx8110, nx8120, nx8134, 
      nx8144, nx8148, booth_integrtaion_1_booth_output_23, nx2991, nx8158, 
      nx8168, nx8182, nx8192, nx8196, booth_integrtaion_1_booth_output_25, 
      nx2993, nx8206, nx8216, nx8230, nx8240, nx8244, 
      booth_integrtaion_1_booth_output_27, nx2995, nx8254, nx8264, nx8278, 
      nx8288, nx8292, booth_integrtaion_1_booth_output_29, nx2997, nx8302, 
      nx8312, booth_integrtaion_1_booth_output_31, nx8326, nx8336, nx8340, 
      nx8342, nx8350, nx8356, nx8368, nx8376, nx8392, nx8400, nx8416, nx8424, 
      nx8440, nx8448, nx8464, nx8472, nx8488, nx8496, nx8508, nx8524, nx8530, 
      nx8536, nx8554, nx8566, nx8578, nx8590, nx8602, nx8614, nx8626, nx8638, 
      nx8650, nx8662, nx8674, nx8686, nx8698, nx8710, nx8722, nx8730, nx8744, 
      nx8746, nx8760, nx8762, nx8776, nx8778, nx8792, nx8794, nx8808, nx8810, 
      nx8824, nx8826, nx8840, booth_integration_output_0_0, 
      booth_integrtaion_0_shift_reg_output_9, 
      booth_integrtaion_0_shift_Reg_count_9, 
      booth_integrtaion_0_shift_Reg_output_8, 
      booth_integrtaion_0_shift_Reg_count_8, 
      booth_integrtaion_0_shift_Reg_output_7, 
      booth_integrtaion_0_shift_Reg_count_7, 
      booth_integrtaion_0_shift_Reg_output_6, 
      booth_integrtaion_0_shift_Reg_count_6, 
      booth_integrtaion_0_shift_Reg_output_5, 
      booth_integrtaion_0_shift_Reg_count_5, 
      booth_integrtaion_0_shift_Reg_output_4, 
      booth_integrtaion_0_shift_Reg_count_4, 
      booth_integrtaion_0_shift_Reg_output_3, 
      booth_integrtaion_0_shift_Reg_count_3, 
      booth_integrtaion_0_shift_Reg_output_2, 
      booth_integrtaion_0_shift_Reg_count_2, 
      booth_integrtaion_0_shift_Reg_output_1, 
      booth_integrtaion_0_shift_Reg_count_1, 
      booth_integrtaion_0_shift_reg_output_0, 
      booth_integrtaion_0_shift_Reg_count_0, booth_integration_output_0_1, 
      booth_integration_output_0_2, booth_integration_output_0_3, 
      booth_integration_output_0_4, booth_integration_output_0_5, 
      booth_integration_output_0_6, booth_integration_output_0_7, 
      booth_integration_output_0_8, booth_integration_output_0_9, 
      booth_integration_output_0_10, booth_integration_output_0_11, 
      booth_integration_output_0_12, booth_integration_output_0_13, 
      booth_integration_output_0_14, booth_integration_output_0_15, 
      booth_integrtaion_0_booth_output_16, nx8976, nx8980, nx8986, 
      booth_integrtaion_0_booth_output_17, nx3000, nx8994, nx9010, nx3001, 
      nx9020, nx9024, nx9038, booth_integrtaion_0_booth_output_19, nx3002, 
      nx9048, nx9058, nx9072, nx9082, nx9086, 
      booth_integrtaion_0_booth_output_21, nx3004, nx9096, nx9106, nx9120, 
      nx9130, nx9134, booth_integrtaion_0_booth_output_23, nx3006, nx9144, 
      nx9154, nx9168, nx9178, nx9182, booth_integrtaion_0_booth_output_25, 
      nx3008, nx9192, nx9202, nx9216, nx9226, nx9230, 
      booth_integrtaion_0_booth_output_27, nx3010, nx9240, nx9250, nx9264, 
      nx9274, nx9278, booth_integrtaion_0_booth_output_29, nx3012, nx9288, 
      nx9298, booth_integrtaion_0_booth_output_31, nx9312, nx9322, nx9326, 
      nx9328, nx9336, nx9342, nx9354, nx9362, nx9378, nx9386, nx9402, nx9410, 
      nx9426, nx9434, nx9450, nx9458, nx9474, nx9482, nx9494, nx9510, nx9516, 
      nx9522, nx9540, nx9552, nx9564, nx9576, nx9588, nx9600, nx9612, nx9624, 
      nx9636, nx9648, nx9660, nx9672, nx9684, nx9696, nx9708, nx9716, nx9730, 
      nx9732, nx9746, nx9748, nx9762, nx9764, nx9778, nx9780, nx9794, nx9796, 
      nx9810, nx9812, nx9826, shift_Reg_adder_0_output_17, 
      shift_Reg_adder_0_output_16, shift_Reg_adder_0_output_15, 
      shift_Reg_adder_0_output_14, shift_Reg_adder_0_output_13, 
      shift_Reg_adder_0_output_12, shift_Reg_adder_0_output_11, 
      shift_Reg_adder_0_output_10, shift_Reg_adder_0_output_9, 
      shift_Reg_adder_0_output_8, shift_Reg_adder_0_output_7, 
      shift_Reg_adder_0_output_6, shift_Reg_adder_0_output_5, 
      shift_Reg_adder_0_output_4, shift_Reg_adder_0_output_3, 
      shift_Reg_adder_0_output_2, shift_Reg_adder_0_output_1, 
      shift_Reg_adder_0_output_0, nx3021, nx3027, nx3041, nx3051, nx3061, 
      nx3071, nx3081, nx3091, nx3101, nx3111, nx3121, nx3131, nx3141, nx3151, 
      nx3161, nx3171, nx3181, nx3191, nx3201, nx3211, nx3221, nx3231, nx3241, 
      nx3251, nx3261, nx3271, nx3281, nx3291, nx3301, nx3311, nx3321, nx3331, 
      nx3341, nx3351, nx3361, nx3371, nx3381, nx3391, nx3401, nx3411, nx3421, 
      nx3431, nx3441, nx3451, nx3461, nx3471, nx3481, nx3491, nx3501, nx3511, 
      nx3521, nx3531, nx3541, nx3551, nx3557, nx3571, nx3581, nx3591, nx3601, 
      nx3611, nx3621, nx3631, nx3641, nx3651, nx3661, nx3671, nx3681, nx3691, 
      nx3701, nx3711, nx3721, nx3731, nx3741, nx3751, nx3761, nx3771, nx3781, 
      nx3791, nx3801, nx3811, nx3821, nx3831, nx3841, nx3851, nx3861, nx3871, 
      nx3881, nx3891, nx3901, nx3911, nx3921, nx3931, nx3941, nx3951, nx3961, 
      nx3971, nx3981, nx3991, nx4001, nx4011, nx4021, nx4031, nx4041, nx4051, 
      nx4061, nx4071, nx4081, nx4087, nx4101, nx4111, nx4121, nx4131, nx4141, 
      nx4151, nx4161, nx4171, nx4181, nx4191, nx4201, nx4211, nx4221, nx4231, 
      nx4241, nx4251, nx4261, nx4271, nx4281, nx4291, nx4301, nx4311, nx4321, 
      nx4331, nx4341, nx4351, nx4361, nx4371, nx4381, nx4391, nx4401, nx4411, 
      nx4421, nx4431, nx4441, nx4451, nx4461, nx4471, nx4481, nx4491, nx4501, 
      nx4511, nx4521, nx4531, nx4541, nx4551, nx4561, nx4571, nx4581, nx4591, 
      nx4601, nx4611, nx4617, nx4631, nx4641, nx4651, nx4661, nx4671, nx4681, 
      nx4691, nx4701, nx4711, nx4721, nx4731, nx4741, nx4751, nx4761, nx4771, 
      nx4781, nx4791, nx4801, nx4811, nx4821, nx4831, nx4841, nx4851, nx4861, 
      nx4871, nx4881, nx4891, nx4901, nx4911, nx4921, nx4931, nx4941, nx4951, 
      nx4961, nx4971, nx4981, nx4991, nx5001, nx5011, nx5021, nx5031, nx5041, 
      nx5051, nx5061, nx5071, nx5081, nx5091, nx5101, nx5111, nx5121, nx5131, 
      nx5141, nx5147, nx5161, nx5171, nx5181, nx5191, nx5201, nx5211, nx5221, 
      nx5231, nx5241, nx5251, nx5261, nx5271, nx5281, nx5291, nx5301, nx5311, 
      nx5321, nx5331, nx5341, nx5351, nx5361, nx5371, nx5381, nx5391, nx5401, 
      nx5411, nx5421, nx5431, nx5441, nx5451, nx5461, nx5471, nx5481, nx5491, 
      nx5501, nx5511, nx5521, nx5531, nx5541, nx5551, nx5561, nx5571, nx5581, 
      nx5591, nx5601, nx5611, nx5621, nx5631, nx5641, nx5651, nx5661, nx5671, 
      nx5677, nx5691, nx5701, nx5711, nx5721, nx5731, nx5741, nx5751, nx5761, 
      nx5771, nx5781, nx5791, nx5801, nx5811, nx5821, nx5831, nx5841, nx5851, 
      nx5861, nx5871, nx5881, nx5891, nx5901, nx5911, nx5921, nx5931, nx5941, 
      nx5951, nx5961, nx5971, nx5981, nx5991, nx6001, nx6011, nx6021, nx6031, 
      nx6041, nx6051, nx6061, nx6071, nx6081, nx6091, nx6101, nx6111, nx6121, 
      nx6131, nx6141, nx6151, nx6161, nx6171, nx6181, nx6191, nx6201, nx6207, 
      nx6221, nx6231, nx6241, nx6251, nx6261, nx6271, nx6281, nx6291, nx6301, 
      nx6311, nx6321, nx6331, nx6341, nx6351, nx6361, nx6371, nx6381, nx6391, 
      nx6401, nx6411, nx6421, nx6431, nx6441, nx6451, nx6461, nx6471, nx6481, 
      nx6491, nx6501, nx6511, nx6521, nx6531, nx6541, nx6551, nx6561, nx6571, 
      nx6581, nx6591, nx6601, nx6611, nx6621, nx6631, nx6641, nx6651, nx6661, 
      nx6671, nx6681, nx6691, nx6701, nx6711, nx6721, nx6731, nx6737, nx6751, 
      nx6761, nx6771, nx6781, nx6791, nx6801, nx6811, nx6821, nx6831, nx6841, 
      nx6851, nx6861, nx6871, nx6881, nx6891, nx6901, nx6911, nx6921, nx6931, 
      nx6941, nx6951, nx6961, nx6971, nx6981, nx6991, nx7001, nx7011, nx7021, 
      nx7031, nx7041, nx7051, nx7061, nx7071, nx7081, nx7091, nx7101, nx7111, 
      nx7121, nx7131, nx7141, nx7151, nx7161, nx7171, nx7181, nx7191, nx7201, 
      nx7211, nx7221, nx7231, nx7241, nx7251, nx7261, nx7267, nx7281, nx7291, 
      nx7301, nx7311, nx7321, nx7331, nx7341, nx7351, nx7361, nx7371, nx7381, 
      nx7391, nx7401, nx7411, nx7421, nx7431, nx7441, nx7451, nx7461, nx7471, 
      nx7481, nx7491, nx7501, nx7511, nx7521, nx7531, nx7541, nx7551, nx7561, 
      nx7571, nx7581, nx7591, nx7601, nx7611, nx7621, nx7631, nx7641, nx7651, 
      nx7661, nx7671, nx7681, nx7691, nx7701, nx7711, nx7721, nx7731, nx7741, 
      nx7751, nx7761, nx7771, nx7781, nx7791, nx7797, nx7811, nx7821, nx7831, 
      nx7841, nx7851, nx7861, nx7871, nx7881, nx7891, nx7901, nx7911, nx7921, 
      nx7931, nx7941, nx7951, nx7961, nx7971, nx7981, nx7991, nx8001, nx8011, 
      nx8021, nx8031, nx8041, nx8051, nx8061, nx8071, nx8081, nx8091, nx8101, 
      nx8111, nx8121, nx8131, nx8141, nx8151, nx8161, nx8171, nx8181, nx8191, 
      nx8201, nx8211, nx8221, nx8231, nx8241, nx8251, nx8261, nx8271, nx8281, 
      nx8291, nx8301, nx8311, done_EXMPLR, nx8321, nx8327, nx8341, nx8351, 
      nx8361, nx8371, nx8381, nx8391, nx8401, nx8411, nx8421, nx8431, nx8441, 
      nx8451, nx8461, nx8471, nx8481, nx8491, nx8501, nx8511, nx8605, nx8668, 
      nx8731, nx8769, nx8777, nx8779, nx8785, nx8791, nx8801, nx8803, nx8807, 
      nx8813, nx8821, nx8823, nx8829, nx8831, nx8835, nx8837, nx8845, nx8847, 
      nx8851, nx8859, nx8865, nx8871, nx8873, nx8879, nx8886, nx8888, nx8893, 
      nx8895, nx8898, nx8902, nx8905, nx8909, nx8911, nx8915, nx8922, nx8924, 
      nx8929, nx8931, nx8934, nx8938, nx8941, nx8945, nx8947, nx8951, nx8958, 
      nx8960, nx8965, nx8967, nx8971, nx8975, nx8979, nx8985, nx8987, nx8993, 
      nx9001, nx9003, nx9011, nx9013, nx9017, nx9023, nx9027, nx9033, nx9035, 
      nx9041, nx9049, nx9051, nx9059, nx9061, nx9065, nx9071, nx9075, nx9083, 
      nx9087, nx9089, nx9097, nx9101, nx9109, nx9113, nx9117, nx9121, nx9125, 
      nx9129, nx9133, nx9139, nx9141, nx9143, nx9146, nx9149, nx9153, nx9157, 
      nx9161, nx9165, nx9167, nx9171, nx9175, nx9181, nx9183, nx9187, nx9191, 
      nx9197, nx9199, nx9203, nx9207, nx9213, nx9215, nx9219, nx9223, nx9229, 
      nx9231, nx9235, nx9239, nx9245, nx9247, nx9251, nx9255, nx9261, nx9263, 
      nx9267, nx9271, nx9277, nx9279, nx9283, nx9361, nx9423, nx9447, nx9453, 
      nx9455, nx9461, nx9466, nx9475, nx9477, nx9480, nx9487, nx9492, nx9495, 
      nx9499, nx9501, nx9504, nx9507, nx9513, nx9515, nx9519, nx9527, nx9532, 
      nx9537, nx9539, nx9544, nx9551, nx9553, nx9558, nx9561, nx9565, nx9569, 
      nx9573, nx9579, nx9581, nx9585, nx9593, nx9595, nx9603, nx9605, nx9609, 
      nx9615, nx9618, nx9623, nx9625, nx9629, nx9637, nx9639, nx9645, nx9647, 
      nx9651, nx9655, nx9659, nx9664, nx9666, nx9671, nx9679, nx9681, nx9688, 
      nx9690, nx9693, nx9699, nx9702, nx9707, nx9709, nx9713, nx9721, nx9723, 
      nx9731, nx9733, nx9737, nx9743, nx9747, nx9755, nx9759, nx9761, nx9769, 
      nx9773, nx9781, nx9785, nx9789, nx9793, nx9797, nx9801, nx9805, nx9811, 
      nx9813, nx9817, nx9821, nx9825, nx9829, nx9831, nx9833, nx9837, nx9839, 
      nx9843, nx9847, nx9853, nx9855, nx9859, nx9863, nx9868, nx9870, nx9874, 
      nx9877, nx9881, nx9883, nx9886, nx9889, nx9893, nx9895, nx9898, nx9901, 
      nx9905, nx9907, nx9910, nx9913, nx9917, nx9919, nx9922, nx9925, nx9929, 
      nx9931, nx9934, nx9982, nx10029, nx10050, nx10055, nx10057, nx10061, 
      nx10065, nx10071, nx10073, nx10076, nx10080, nx10085, nx10087, nx10091, 
      nx10093, nx10096, nx10098, nx10103, nx10105, nx10108, nx10114, nx10119, 
      nx10123, nx10125, nx10129, nx10136, nx10138, nx10143, nx10145, nx10148, 
      nx10152, nx10155, nx10159, nx10161, nx10165, nx10172, nx10174, nx10179, 
      nx10181, nx10184, nx10188, nx10191, nx10195, nx10197, nx10201, nx10208, 
      nx10210, nx10215, nx10217, nx10220, nx10224, nx10227, nx10231, nx10233, 
      nx10237, nx10244, nx10246, nx10251, nx10253, nx10256, nx10260, nx10263, 
      nx10267, nx10269, nx10273, nx10280, nx10282, nx10287, nx10289, nx10292, 
      nx10296, nx10299, nx10304, nx10307, nx10309, nx10316, nx10319, nx10324, 
      nx10328, nx10332, nx10336, nx10340, nx10344, nx10347, nx10351, nx10353, 
      nx10355, nx10357, nx10359, nx10361, nx10363, nx10365, nx10368, nx10370, 
      nx10373, nx10376, nx10380, nx10382, nx10385, nx10388, nx10392, nx10394, 
      nx10397, nx10400, nx10404, nx10406, nx10409, nx10412, nx10416, nx10418, 
      nx10421, nx10424, nx10428, nx10430, nx10433, nx10436, nx10440, nx10442, 
      nx10445, nx10448, nx10452, nx10454, nx10457, nx10505, nx10552, nx10573, 
      nx10578, nx10580, nx10584, nx10588, nx10594, nx10596, nx10599, nx10603, 
      nx10608, nx10610, nx10614, nx10616, nx10619, nx10621, nx10626, nx10628, 
      nx10631, nx10637, nx10642, nx10646, nx10648, nx10652, nx10659, nx10661, 
      nx10666, nx10668, nx10671, nx10675, nx10678, nx10682, nx10684, nx10688, 
      nx10695, nx10697, nx10702, nx10704, nx10707, nx10711, nx10714, nx10718, 
      nx10720, nx10724, nx10731, nx10733, nx10738, nx10740, nx10743, nx10747, 
      nx10750, nx10754, nx10756, nx10760, nx10767, nx10769, nx10774, nx10776, 
      nx10779, nx10783, nx10786, nx10790, nx10792, nx10796, nx10803, nx10805, 
      nx10810, nx10812, nx10815, nx10819, nx10822, nx10827, nx10830, nx10832, 
      nx10839, nx10842, nx10847, nx10851, nx10855, nx10859, nx10863, nx10867, 
      nx10870, nx10874, nx10876, nx10878, nx10880, nx10882, nx10884, nx10886, 
      nx10888, nx10891, nx10893, nx10896, nx10899, nx10903, nx10905, nx10908, 
      nx10911, nx10915, nx10917, nx10920, nx10923, nx10927, nx10929, nx10932, 
      nx10935, nx10939, nx10941, nx10944, nx10947, nx10951, nx10953, nx10956, 
      nx10959, nx10963, nx10965, nx10968, nx10971, nx10975, nx10977, nx10980, 
      nx11028, nx11075, nx11096, nx11101, nx11103, nx11107, nx11111, nx11117, 
      nx11119, nx11122, nx11126, nx11131, nx11133, nx11137, nx11139, nx11142, 
      nx11144, nx11149, nx11151, nx11154, nx11160, nx11165, nx11169, nx11171, 
      nx11175, nx11182, nx11184, nx11189, nx11191, nx11194, nx11198, nx11201, 
      nx11205, nx11207, nx11211, nx11218, nx11220, nx11225, nx11227, nx11230, 
      nx11234, nx11237, nx11241, nx11243, nx11247, nx11254, nx11256, nx11261, 
      nx11263, nx11266, nx11270, nx11273, nx11277, nx11279, nx11283, nx11290, 
      nx11292, nx11297, nx11299, nx11302, nx11306, nx11309, nx11313, nx11315, 
      nx11319, nx11326, nx11328, nx11333, nx11335, nx11338, nx11342, nx11345, 
      nx11350, nx11353, nx11355, nx11362, nx11365, nx11370, nx11374, nx11378, 
      nx11382, nx11386, nx11390, nx11393, nx11397, nx11399, nx11401, nx11403, 
      nx11405, nx11407, nx11409, nx11411, nx11414, nx11416, nx11419, nx11422, 
      nx11426, nx11428, nx11431, nx11434, nx11438, nx11440, nx11443, nx11446, 
      nx11450, nx11452, nx11455, nx11458, nx11462, nx11464, nx11467, nx11470, 
      nx11474, nx11476, nx11479, nx11482, nx11486, nx11488, nx11491, nx11494, 
      nx11498, nx11500, nx11503, nx11551, nx11598, nx11619, nx11624, nx11626, 
      nx11630, nx11634, nx11640, nx11642, nx11645, nx11649, nx11654, nx11656, 
      nx11660, nx11662, nx11665, nx11667, nx11672, nx11674, nx11677, nx11683, 
      nx11688, nx11692, nx11694, nx11698, nx11705, nx11707, nx11712, nx11714, 
      nx11717, nx11721, nx11724, nx11728, nx11730, nx11734, nx11741, nx11743, 
      nx11748, nx11750, nx11753, nx11757, nx11760, nx11764, nx11766, nx11770, 
      nx11777, nx11779, nx11784, nx11786, nx11789, nx11793, nx11796, nx11800, 
      nx11802, nx11806, nx11813, nx11815, nx11820, nx11822, nx11825, nx11829, 
      nx11832, nx11836, nx11838, nx11842, nx11849, nx11851, nx11856, nx11858, 
      nx11861, nx11865, nx11868, nx11873, nx11876, nx11878, nx11885, nx11888, 
      nx11893, nx11897, nx11901, nx11905, nx11909, nx11913, nx11916, nx11920, 
      nx11922, nx11924, nx11926, nx11928, nx11930, nx11932, nx11934, nx11937, 
      nx11939, nx11942, nx11945, nx11949, nx11951, nx11954, nx11957, nx11961, 
      nx11963, nx11966, nx11969, nx11973, nx11975, nx11978, nx11981, nx11985, 
      nx11987, nx11990, nx11993, nx11997, nx11999, nx12002, nx12005, nx12009, 
      nx12011, nx12014, nx12017, nx12021, nx12023, nx12026, nx12074, nx12121, 
      nx12142, nx12147, nx12149, nx12153, nx12157, nx12163, nx12165, nx12168, 
      nx12172, nx12177, nx12179, nx12183, nx12185, nx12188, nx12190, nx12195, 
      nx12197, nx12200, nx12206, nx12211, nx12215, nx12217, nx12221, nx12228, 
      nx12230, nx12235, nx12237, nx12240, nx12244, nx12247, nx12251, nx12253, 
      nx12257, nx12264, nx12266, nx12271, nx12273, nx12276, nx12280, nx12283, 
      nx12287, nx12289, nx12293, nx12300, nx12302, nx12307, nx12309, nx12312, 
      nx12316, nx12319, nx12323, nx12325, nx12329, nx12336, nx12338, nx12343, 
      nx12345, nx12348, nx12352, nx12355, nx12359, nx12361, nx12365, nx12372, 
      nx12374, nx12379, nx12381, nx12384, nx12388, nx12391, nx12396, nx12399, 
      nx12401, nx12408, nx12411, nx12416, nx12420, nx12424, nx12428, nx12432, 
      nx12436, nx12439, nx12443, nx12445, nx12447, nx12449, nx12451, nx12453, 
      nx12455, nx12457, nx12460, nx12462, nx12465, nx12468, nx12472, nx12474, 
      nx12477, nx12480, nx12484, nx12486, nx12489, nx12492, nx12496, nx12498, 
      nx12501, nx12504, nx12508, nx12510, nx12513, nx12516, nx12520, nx12522, 
      nx12525, nx12528, nx12532, nx12534, nx12537, nx12540, nx12544, nx12546, 
      nx12549, nx12597, nx12644, nx12665, nx12670, nx12672, nx12676, nx12680, 
      nx12686, nx12688, nx12691, nx12695, nx12700, nx12702, nx12706, nx12708, 
      nx12711, nx12713, nx12718, nx12720, nx12723, nx12729, nx12734, nx12738, 
      nx12740, nx12744, nx12751, nx12753, nx12758, nx12760, nx12763, nx12767, 
      nx12770, nx12774, nx12776, nx12780, nx12787, nx12789, nx12794, nx12796, 
      nx12799, nx12803, nx12806, nx12810, nx12812, nx12816, nx12823, nx12825, 
      nx12830, nx12832, nx12835, nx12839, nx12842, nx12846, nx12848, nx12852, 
      nx12859, nx12861, nx12866, nx12868, nx12871, nx12875, nx12878, nx12882, 
      nx12884, nx12888, nx12895, nx12897, nx12902, nx12904, nx12907, nx12911, 
      nx12914, nx12919, nx12922, nx12924, nx12931, nx12934, nx12939, nx12943, 
      nx12947, nx12951, nx12955, nx12959, nx12962, nx12966, nx12968, nx12970, 
      nx12972, nx12974, nx12976, nx12978, nx12980, nx12983, nx12985, nx12988, 
      nx12991, nx12995, nx12997, nx13000, nx13003, nx13007, nx13009, nx13012, 
      nx13015, nx13019, nx13021, nx13024, nx13027, nx13031, nx13033, nx13036, 
      nx13039, nx13043, nx13045, nx13048, nx13051, nx13055, nx13057, nx13060, 
      nx13063, nx13067, nx13069, nx13072, nx13120, nx13167, nx13188, nx13193, 
      nx13195, nx13199, nx13203, nx13209, nx13211, nx13214, nx13218, nx13223, 
      nx13225, nx13229, nx13231, nx13234, nx13236, nx13241, nx13243, nx13246, 
      nx13252, nx13257, nx13261, nx13263, nx13267, nx13274, nx13276, nx13281, 
      nx13283, nx13286, nx13290, nx13293, nx13297, nx13299, nx13303, nx13310, 
      nx13312, nx13317, nx13319, nx13322, nx13326, nx13329, nx13333, nx13335, 
      nx13339, nx13346, nx13348, nx13353, nx13355, nx13358, nx13362, nx13365, 
      nx13369, nx13371, nx13375, nx13382, nx13384, nx13389, nx13391, nx13394, 
      nx13398, nx13401, nx13405, nx13407, nx13411, nx13418, nx13420, nx13425, 
      nx13427, nx13430, nx13434, nx13437, nx13442, nx13445, nx13447, nx13454, 
      nx13457, nx13462, nx13466, nx13470, nx13474, nx13478, nx13482, nx13485, 
      nx13489, nx13491, nx13493, nx13495, nx13497, nx13499, nx13501, nx13503, 
      nx13506, nx13508, nx13511, nx13514, nx13518, nx13520, nx13523, nx13526, 
      nx13530, nx13532, nx13535, nx13538, nx13542, nx13544, nx13547, nx13550, 
      nx13554, nx13556, nx13559, nx13562, nx13566, nx13568, nx13571, nx13574, 
      nx13578, nx13580, nx13583, nx13586, nx13590, nx13592, nx13595, nx13643, 
      nx13690, nx13711, nx13716, nx13718, nx13722, nx13726, nx13732, nx13734, 
      nx13737, nx13741, nx13746, nx13748, nx13752, nx13754, nx13757, nx13759, 
      nx13764, nx13766, nx13769, nx13775, nx13780, nx13784, nx13786, nx13790, 
      nx13797, nx13799, nx13804, nx13806, nx13809, nx13813, nx13816, nx13820, 
      nx13822, nx13826, nx13833, nx13835, nx13840, nx13842, nx13845, nx13849, 
      nx13852, nx13856, nx13858, nx13862, nx13869, nx13871, nx13876, nx13878, 
      nx13881, nx13885, nx13888, nx13892, nx13894, nx13898, nx13905, nx13907, 
      nx13912, nx13914, nx13917, nx13921, nx13924, nx13928, nx13930, nx13934, 
      nx13941, nx13943, nx13948, nx13950, nx13953, nx13957, nx13960, nx13965, 
      nx13968, nx13970, nx13977, nx13980, nx13985, nx13989, nx13993, nx13997, 
      nx14001, nx14005, nx14008, nx14012, nx14014, nx14016, nx14018, nx14020, 
      nx14022, nx14024, nx14026, nx14029, nx14031, nx14034, nx14037, nx14041, 
      nx14043, nx14046, nx14049, nx14053, nx14055, nx14058, nx14061, nx14065, 
      nx14067, nx14070, nx14073, nx14077, nx14079, nx14082, nx14085, nx14089, 
      nx14091, nx14094, nx14097, nx14101, nx14103, nx14106, nx14109, nx14113, 
      nx14115, nx14122, nx14136, nx14138, nx14140, nx14142, nx14144, nx14146, 
      nx14148, nx14150, nx14152, nx14154, nx14156, nx14158, nx14160, nx14162, 
      nx14164, nx14166, nx14168, nx14170, nx14172, nx14174, nx14182, nx14196, 
      nx14204, nx14218, nx14226, nx14240, nx14248, nx14262, nx14270, nx14284, 
      nx14292, nx14306, nx14314, nx14328, nx14336, nx14350, nx14358, nx14372, 
      nx14382, nx14388, nx14390, nx14392, nx14394, nx14396, nx14400, nx14402, 
      nx14404, nx14406, nx14408, nx14410, nx14412, nx14414, nx14416, nx14418, 
      nx14422, nx14424, nx14426, nx14428, nx14430, nx14432, nx14434, nx14436, 
      nx14438, nx14440, nx14444, nx14446, nx14448, nx14450, nx14452, nx14454, 
      nx14456, nx14458, nx14460, nx14462, nx14466, nx14468, nx14470, nx14472, 
      nx14474, nx14476, nx14478, nx14480, nx14482, nx14484, nx14488, nx14490, 
      nx14492, nx14494, nx14496, nx14498, nx14500, nx14502, nx14504, nx14506, 
      nx14510, nx14512, nx14514, nx14516, nx14518, nx14520, nx14522, nx14524, 
      nx14526, nx14528, nx14532, nx14534, nx14536, nx14538, nx14540, nx14542, 
      nx14544, nx14546, nx14548, nx14550, nx14554, nx14556, nx14558, nx14560, 
      nx14562, nx14564, nx14566, nx14568, nx14570, nx14572, nx14576, nx14578, 
      nx14580, nx14582, nx14584, nx14586, nx14588, nx14590, nx14592, nx14594, 
      nx14598, nx14600, nx14602, nx14604, nx14606, nx14612, nx14614, nx14616, 
      nx14618, nx14620, nx14622, nx14624, nx14626, nx14628, nx14630, nx14632, 
      nx14634, nx14636, nx14638, nx14640, nx14642, nx14644, nx14646, nx14648, 
      nx14650, nx14652, nx14654, nx14656, nx14658, nx14660, nx14662, nx14664, 
      nx14666, nx14668, nx14670, nx14672, nx14674, nx14676, nx14678, nx14680, 
      nx14682, nx14684, nx14686, nx14688, nx14690, nx14692, nx14694, nx14696, 
      nx14698, nx14700, nx14702, nx14704, nx14706, nx14708, nx14710, nx14712, 
      nx14714, nx14716, nx14718, nx14720, nx14722, nx14724, nx14726, nx14728, 
      nx14730, nx14732, nx14734, nx14736, nx14738, nx14740, nx14742, nx14744, 
      nx14746, nx14748, nx14750, nx14752, nx14754, nx14756, nx14758, nx14760, 
      nx14762, nx14764, nx14766, nx14768, nx14770, nx14772, nx14774, nx14776, 
      nx14778, nx14780, nx14782, nx14784, nx14786, nx14788, nx14790, nx14792, 
      nx14794, nx14796, nx14798, nx14800, nx14802, nx14804, nx14806, nx14808, 
      nx14810, nx14812, nx14814, nx14816, nx14822, nx14824, nx14826, nx14828, 
      nx14830, nx14832, nx14834, nx14836, nx14838, nx14840, nx14842, nx14844, 
      nx14846, nx14848, nx14850, nx14852, nx14854, nx14856, nx14858, nx14860
   : std_logic ;

begin
   done <= done_EXMPLR ;
   dec_enable <= dec_sel_0_EXMPLR ;
   dec_sel(3) <= dec_sel_0_EXMPLR ;
   dec_sel(2) <= dec_sel_0_EXMPLR ;
   dec_sel(1) <= dec_sel_0_EXMPLR ;
   dec_sel(0) <= dec_sel_0_EXMPLR ;
   shift_Reg_adder_0_reg_count_19 : dffr port map ( Q=>done_EXMPLR, QB=>OPEN, 
      D=>nx8321, CLK=>clk, R=>nx14140);
   ix8322 : or02 port map ( Y=>nx8321, A0=>nx14382, A1=>dec_sel_0_EXMPLR);
   shift_Reg_adder_0_reg_count_18 : dffr port map ( Q=>dec_sel_0_EXMPLR, QB
      =>OPEN, D=>nx8511, CLK=>clk, R=>nx14140);
   shift_Reg_adder_0_reg_count_17 : dffr port map ( Q=>
      shift_Reg_adder_0_output_17, QB=>OPEN, D=>nx8501, CLK=>clk, R=>nx14140
   );
   shift_Reg_adder_0_reg_count_16 : dffr port map ( Q=>
      shift_Reg_adder_0_output_16, QB=>OPEN, D=>nx8491, CLK=>clk, R=>nx14140
   );
   shift_Reg_adder_0_reg_count_15 : dffr port map ( Q=>
      shift_Reg_adder_0_output_15, QB=>OPEN, D=>nx8481, CLK=>clk, R=>nx14140
   );
   shift_Reg_adder_0_reg_count_14 : dffr port map ( Q=>
      shift_Reg_adder_0_output_14, QB=>OPEN, D=>nx8471, CLK=>clk, R=>nx14140
   );
   shift_Reg_adder_0_reg_count_13 : dffr port map ( Q=>
      shift_Reg_adder_0_output_13, QB=>OPEN, D=>nx8461, CLK=>clk, R=>nx14138
   );
   shift_Reg_adder_0_reg_count_12 : dffr port map ( Q=>
      shift_Reg_adder_0_output_12, QB=>OPEN, D=>nx8451, CLK=>clk, R=>nx14138
   );
   shift_Reg_adder_0_reg_count_11 : dffr port map ( Q=>
      shift_Reg_adder_0_output_11, QB=>OPEN, D=>nx8441, CLK=>clk, R=>nx14138
   );
   shift_Reg_adder_0_reg_count_10 : dffr port map ( Q=>
      shift_Reg_adder_0_output_10, QB=>OPEN, D=>nx8431, CLK=>clk, R=>nx14138
   );
   shift_Reg_adder_0_reg_count_9 : dffr port map ( Q=>
      shift_Reg_adder_0_output_9, QB=>OPEN, D=>nx8421, CLK=>clk, R=>nx14138
   );
   shift_Reg_adder_0_reg_count_8 : dffr port map ( Q=>
      shift_Reg_adder_0_output_8, QB=>OPEN, D=>nx8411, CLK=>clk, R=>nx14138
   );
   shift_Reg_adder_0_reg_count_7 : dffr port map ( Q=>
      shift_Reg_adder_0_output_7, QB=>OPEN, D=>nx8401, CLK=>clk, R=>nx14138
   );
   shift_Reg_adder_0_reg_count_6 : dffr port map ( Q=>
      shift_Reg_adder_0_output_6, QB=>OPEN, D=>nx8391, CLK=>clk, R=>nx14136
   );
   shift_Reg_adder_0_reg_count_5 : dffr port map ( Q=>
      shift_Reg_adder_0_output_5, QB=>OPEN, D=>nx8381, CLK=>clk, R=>nx14136
   );
   shift_Reg_adder_0_reg_count_4 : dffr port map ( Q=>
      shift_Reg_adder_0_output_4, QB=>OPEN, D=>nx8371, CLK=>clk, R=>nx14136
   );
   shift_Reg_adder_0_reg_count_3 : dffr port map ( Q=>
      shift_Reg_adder_0_output_3, QB=>OPEN, D=>nx8361, CLK=>clk, R=>nx14136
   );
   shift_Reg_adder_0_reg_count_2 : dffr port map ( Q=>
      shift_Reg_adder_0_output_2, QB=>OPEN, D=>nx8351, CLK=>clk, R=>nx14136
   );
   shift_Reg_adder_0_reg_count_1 : dffr port map ( Q=>
      shift_Reg_adder_0_output_1, QB=>OPEN, D=>nx8341, CLK=>clk, R=>nx14136
   );
   shift_Reg_adder_0_reg_count_0 : dffs_ni port map ( Q=>
      shift_Reg_adder_0_output_0, QB=>OPEN, D=>nx8327, CLK=>clk, S=>nx14136
   );
   booth_integrtaion_9_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_1, QB=>OPEN, D=>nx3531, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_2, QB=>nx9161, D=>nx3521, CLK=>clk, R=>rst
   );
   booth_integrtaion_9_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_3, QB=>OPEN, D=>nx3511, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_4, QB=>nx9157, D=>nx3501, CLK=>clk, R=>rst
   );
   booth_integrtaion_9_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_5, QB=>OPEN, D=>nx3491, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_6, QB=>nx9153, D=>nx3481, CLK=>clk, R=>rst
   );
   booth_integrtaion_9_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_7, QB=>OPEN, D=>nx3471, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_8, QB=>nx9149, D=>nx3461, CLK=>clk, R=>rst
   );
   booth_integrtaion_9_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_9, QB=>OPEN, D=>nx3451, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_10, QB=>nx9146, D=>nx3441, CLK=>clk, R=>rst
   );
   booth_integrtaion_9_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_11, QB=>OPEN, D=>nx3431, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_12, QB=>nx9143, D=>nx3421, CLK=>clk, R=>rst
   );
   booth_integrtaion_9_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_13, QB=>OPEN, D=>nx3411, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_14, QB=>nx9141, D=>nx3401, CLK=>clk, R=>rst
   );
   ix8669 : aoi22 port map ( Y=>nx8668, A0=>neuron(15), A1=>nx14174, B0=>
      nx642, B1=>nx648);
   booth_integrtaion_9_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_reg_output_0, QB=>OPEN, D=>nx3041, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_0, QB=>OPEN, D=>nx3027, CLK=>clk, 
      S=>nx14144);
   booth_integrtaion_9_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_reg_output_9, QB=>OPEN, D=>nx3221, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_9, QB=>OPEN, D=>nx3211, CLK=>clk, 
      R=>nx14144);
   booth_integrtaion_9_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_8, QB=>OPEN, D=>nx3201, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_8, QB=>OPEN, D=>nx3191, CLK=>clk, 
      R=>nx14144);
   booth_integrtaion_9_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_7, QB=>OPEN, D=>nx3181, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_7, QB=>OPEN, D=>nx3171, CLK=>clk, 
      R=>nx14142);
   booth_integrtaion_9_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_6, QB=>OPEN, D=>nx3161, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_6, QB=>OPEN, D=>nx3151, CLK=>clk, 
      R=>nx14142);
   booth_integrtaion_9_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_5, QB=>OPEN, D=>nx3141, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_5, QB=>OPEN, D=>nx3131, CLK=>clk, 
      R=>nx14142);
   booth_integrtaion_9_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_4, QB=>OPEN, D=>nx3121, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_4, QB=>OPEN, D=>nx3111, CLK=>clk, 
      R=>nx14142);
   booth_integrtaion_9_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_3, QB=>OPEN, D=>nx3101, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_3, QB=>OPEN, D=>nx3091, CLK=>clk, 
      R=>nx14142);
   booth_integrtaion_9_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_2, QB=>OPEN, D=>nx3081, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_2, QB=>OPEN, D=>nx3071, CLK=>clk, 
      R=>nx14142);
   booth_integrtaion_9_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_output_1, QB=>OPEN, D=>nx3061, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_9_shift_Reg_count_1, QB=>OPEN, D=>nx3051, CLK=>clk, 
      R=>nx14140);
   ix3022 : nand02 port map ( Y=>nx3021, A0=>nx14612, A1=>nx14122);
   booth_integrtaion_9_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx8731, D=>nx3021, CLK=>clk, S=>nx14142);
   ix643 : nand02 port map ( Y=>nx642, A0=>nx8769, A1=>nx8785);
   ix8770 : oai21 port map ( Y=>nx8769, A0=>nx106, A1=>nx102, B0=>
      weight_9(0));
   ix3232 : oai21 port map ( Y=>nx3231, A0=>nx8777, A1=>nx14388, B0=>nx8779
   );
   booth_integrtaion_9_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx8777, D=>nx3231, CLK=>clk, R=>rst);
   booth_integrtaion_9_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_0, QB=>nx8605, D=>nx3541, CLK=>clk, R=>rst
   );
   ix8792 : xnor2 port map ( Y=>nx8791, A0=>nx112, A1=>nx2805);
   ix3372 : oai21 port map ( Y=>nx3371, A0=>nx8801, A1=>nx14388, B0=>nx8803
   );
   booth_integrtaion_9_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_17, QB=>nx8801, D=>nx3371, CLK=>clk, 
      R=>rst);
   ix8804 : nand03 port map ( Y=>nx8803, A0=>nx14396, A1=>nx620, A2=>nx14658
   );
   ix621 : xnor2 port map ( Y=>nx620, A0=>nx8807, A1=>nx2807);
   ix8808 : aoi22 port map ( Y=>nx8807, A0=>
      booth_integrtaion_9_booth_output_17, A1=>nx136, B0=>nx112, B1=>nx2805
   );
   ix121 : nand02 port map ( Y=>nx120, A0=>weight_9(1), A1=>weight_9(0));
   ix8814 : or02 port map ( Y=>nx8813, A0=>weight_9(0), A1=>weight_9(1));
   ix3362 : oai21 port map ( Y=>nx3361, A0=>nx8821, A1=>nx14388, B0=>nx8823
   );
   booth_integrtaion_9_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx8821, D=>nx3361, CLK=>clk, R=>rst);
   ix8824 : nand03 port map ( Y=>nx8823, A0=>nx14396, A1=>nx608, A2=>nx14658
   );
   ix609 : xnor2 port map ( Y=>nx608, A0=>nx164, A1=>nx8837);
   ix165 : oai22 port map ( Y=>nx164, A0=>nx8807, A1=>nx8829, B0=>nx8821, B1
      =>nx14400);
   ix8832 : aoi32 port map ( Y=>nx8831, A0=>nx146, A1=>nx106, A2=>nx8835, B0
      =>weight_9(2), B1=>nx102);
   ix147 : oai21 port map ( Y=>nx146, A0=>weight_9(0), A1=>weight_9(1), B0=>
      weight_9(2));
   ix8838 : xnor2 port map ( Y=>nx8837, A0=>
      booth_integrtaion_9_booth_output_19, A1=>nx184);
   booth_integrtaion_9_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_19, QB=>OPEN, D=>nx3351, CLK=>clk, R
      =>rst);
   ix8846 : xnor2 port map ( Y=>nx8845, A0=>nx8847, A1=>nx8865);
   ix8848 : aoi22 port map ( Y=>nx8847, A0=>
      booth_integrtaion_9_booth_output_19, A1=>nx184, B0=>nx164, B1=>nx2808
   );
   ix185 : oai32 port map ( Y=>nx184, A0=>nx8851, A1=>nx14402, A2=>nx174, B0
      =>nx8859, B1=>nx14406);
   ix8852 : nor02ii port map ( Y=>nx8851, A0=>nx150, A1=>weight_9(3));
   ix151 : nor03_2x port map ( Y=>nx150, A0=>weight_9(2), A1=>weight_9(0), 
      A2=>weight_9(1));
   ix175 : nor04 port map ( Y=>nx174, A0=>weight_9(3), A1=>weight_9(2), A2=>
      weight_9(0), A3=>weight_9(1));
   ix8860 : inv01 port map ( Y=>nx8859, A=>weight_9(3));
   ix3342 : oai21 port map ( Y=>nx3341, A0=>nx8871, A1=>nx14388, B0=>nx8873
   );
   booth_integrtaion_9_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx8871, D=>nx3341, CLK=>clk, R=>rst);
   ix8874 : nand03 port map ( Y=>nx8873, A0=>nx14396, A1=>nx584, A2=>nx14658
   );
   ix585 : xnor2 port map ( Y=>nx584, A0=>nx212, A1=>nx8888);
   ix213 : oai22 port map ( Y=>nx212, A0=>nx8847, A1=>nx8865, B0=>nx8871, B1
      =>nx8879);
   ix8887 : inv01 port map ( Y=>nx8886, A=>weight_9(4));
   ix8889 : xnor2 port map ( Y=>nx8888, A0=>
      booth_integrtaion_9_booth_output_21, A1=>nx232);
   booth_integrtaion_9_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_21, QB=>OPEN, D=>nx3331, CLK=>clk, R
      =>rst);
   ix8894 : xnor2 port map ( Y=>nx8893, A0=>nx8895, A1=>nx8905);
   ix8896 : aoi22 port map ( Y=>nx8895, A0=>
      booth_integrtaion_9_booth_output_21, A1=>nx232, B0=>nx212, B1=>nx2810
   );
   ix233 : oai32 port map ( Y=>nx232, A0=>nx8898, A1=>nx14402, A2=>nx222, B0
      =>nx8902, B1=>nx14406);
   ix8899 : nor02ii port map ( Y=>nx8898, A0=>nx198, A1=>weight_9(5));
   ix199 : nor02ii port map ( Y=>nx198, A0=>weight_9(4), A1=>nx174);
   ix223 : nor02ii port map ( Y=>nx222, A0=>weight_9(5), A1=>nx198);
   ix8903 : inv01 port map ( Y=>nx8902, A=>weight_9(5));
   ix3322 : oai21 port map ( Y=>nx3321, A0=>nx8909, A1=>nx14388, B0=>nx8911
   );
   booth_integrtaion_9_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx8909, D=>nx3321, CLK=>clk, R=>rst);
   ix8912 : nand03 port map ( Y=>nx8911, A0=>nx14396, A1=>nx560, A2=>nx14390
   );
   ix561 : xnor2 port map ( Y=>nx560, A0=>nx260, A1=>nx8924);
   ix261 : oai22 port map ( Y=>nx260, A0=>nx8895, A1=>nx8905, B0=>nx8909, B1
      =>nx8915);
   ix8923 : inv01 port map ( Y=>nx8922, A=>weight_9(6));
   ix8925 : xnor2 port map ( Y=>nx8924, A0=>
      booth_integrtaion_9_booth_output_23, A1=>nx280);
   booth_integrtaion_9_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_23, QB=>OPEN, D=>nx3311, CLK=>clk, R
      =>rst);
   ix8930 : xnor2 port map ( Y=>nx8929, A0=>nx8931, A1=>nx8941);
   ix8932 : aoi22 port map ( Y=>nx8931, A0=>
      booth_integrtaion_9_booth_output_23, A1=>nx280, B0=>nx260, B1=>nx2813
   );
   ix281 : oai32 port map ( Y=>nx280, A0=>nx8934, A1=>nx14402, A2=>nx270, B0
      =>nx8938, B1=>nx14406);
   ix8935 : nor02ii port map ( Y=>nx8934, A0=>nx246, A1=>weight_9(7));
   ix247 : nor02ii port map ( Y=>nx246, A0=>weight_9(6), A1=>nx222);
   ix271 : nor02ii port map ( Y=>nx270, A0=>weight_9(7), A1=>nx246);
   ix8939 : inv01 port map ( Y=>nx8938, A=>weight_9(7));
   ix3302 : oai21 port map ( Y=>nx3301, A0=>nx8945, A1=>nx14390, B0=>nx8947
   );
   booth_integrtaion_9_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx8945, D=>nx3301, CLK=>clk, R=>rst);
   ix8948 : nand03 port map ( Y=>nx8947, A0=>nx14396, A1=>nx536, A2=>nx14390
   );
   ix537 : xnor2 port map ( Y=>nx536, A0=>nx308, A1=>nx8960);
   ix309 : oai22 port map ( Y=>nx308, A0=>nx8931, A1=>nx8941, B0=>nx8945, B1
      =>nx8951);
   ix8959 : inv01 port map ( Y=>nx8958, A=>weight_9(8));
   ix8961 : xnor2 port map ( Y=>nx8960, A0=>
      booth_integrtaion_9_booth_output_25, A1=>nx328);
   booth_integrtaion_9_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_25, QB=>OPEN, D=>nx3291, CLK=>clk, R
      =>rst);
   ix8966 : xnor2 port map ( Y=>nx8965, A0=>nx8967, A1=>nx8979);
   ix8968 : aoi22 port map ( Y=>nx8967, A0=>
      booth_integrtaion_9_booth_output_25, A1=>nx328, B0=>nx308, B1=>nx2817
   );
   ix329 : oai32 port map ( Y=>nx328, A0=>nx8971, A1=>nx14402, A2=>nx318, B0
      =>nx8975, B1=>nx14406);
   ix8972 : nor02ii port map ( Y=>nx8971, A0=>nx294, A1=>weight_9(9));
   ix295 : nor02ii port map ( Y=>nx294, A0=>weight_9(8), A1=>nx270);
   ix319 : nor02ii port map ( Y=>nx318, A0=>weight_9(9), A1=>nx294);
   ix8976 : inv01 port map ( Y=>nx8975, A=>weight_9(9));
   ix3282 : oai21 port map ( Y=>nx3281, A0=>nx8985, A1=>nx14390, B0=>nx8987
   );
   booth_integrtaion_9_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx8985, D=>nx3281, CLK=>clk, R=>rst);
   ix8988 : nand03 port map ( Y=>nx8987, A0=>nx14396, A1=>nx512, A2=>nx14390
   );
   ix513 : xnor2 port map ( Y=>nx512, A0=>nx356, A1=>nx9003);
   ix357 : oai22 port map ( Y=>nx356, A0=>nx8967, A1=>nx8979, B0=>nx8985, B1
      =>nx8993);
   ix9002 : inv01 port map ( Y=>nx9001, A=>weight_9(10));
   ix9004 : xnor2 port map ( Y=>nx9003, A0=>
      booth_integrtaion_9_booth_output_27, A1=>nx376);
   booth_integrtaion_9_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_27, QB=>OPEN, D=>nx3271, CLK=>clk, R
      =>rst);
   ix9012 : xnor2 port map ( Y=>nx9011, A0=>nx9013, A1=>nx9027);
   ix9014 : aoi22 port map ( Y=>nx9013, A0=>
      booth_integrtaion_9_booth_output_27, A1=>nx376, B0=>nx356, B1=>nx2821
   );
   ix377 : oai32 port map ( Y=>nx376, A0=>nx9017, A1=>nx14402, A2=>nx366, B0
      =>nx9023, B1=>nx14406);
   ix9018 : nor02ii port map ( Y=>nx9017, A0=>nx342, A1=>weight_9(11));
   ix343 : nor02ii port map ( Y=>nx342, A0=>weight_9(10), A1=>nx318);
   ix367 : nor02ii port map ( Y=>nx366, A0=>weight_9(11), A1=>nx342);
   ix9024 : inv01 port map ( Y=>nx9023, A=>weight_9(11));
   ix3262 : oai21 port map ( Y=>nx3261, A0=>nx9033, A1=>nx14390, B0=>nx9035
   );
   booth_integrtaion_9_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9033, D=>nx3261, CLK=>clk, R=>rst);
   ix9036 : nand03 port map ( Y=>nx9035, A0=>nx14666, A1=>nx488, A2=>nx14390
   );
   ix489 : xnor2 port map ( Y=>nx488, A0=>nx404, A1=>nx9051);
   ix405 : oai22 port map ( Y=>nx404, A0=>nx9013, A1=>nx9027, B0=>nx9033, B1
      =>nx9041);
   ix9050 : inv01 port map ( Y=>nx9049, A=>weight_9(12));
   ix9052 : xnor2 port map ( Y=>nx9051, A0=>
      booth_integrtaion_9_booth_output_29, A1=>nx424);
   booth_integrtaion_9_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_29, QB=>OPEN, D=>nx3251, CLK=>clk, R
      =>rst);
   ix9060 : xnor2 port map ( Y=>nx9059, A0=>nx9061, A1=>nx9075);
   ix9062 : aoi22 port map ( Y=>nx9061, A0=>
      booth_integrtaion_9_booth_output_29, A1=>nx424, B0=>nx404, B1=>nx2825
   );
   ix425 : oai32 port map ( Y=>nx424, A0=>nx9065, A1=>nx14402, A2=>nx414, B0
      =>nx9071, B1=>nx14406);
   ix9066 : nor02ii port map ( Y=>nx9065, A0=>nx390, A1=>weight_9(13));
   ix391 : nor02ii port map ( Y=>nx390, A0=>weight_9(12), A1=>nx366);
   ix415 : nor02ii port map ( Y=>nx414, A0=>weight_9(13), A1=>nx390);
   ix9072 : inv01 port map ( Y=>nx9071, A=>weight_9(13));
   ix9084 : xnor2 port map ( Y=>nx9083, A0=>nx452, A1=>nx462);
   ix453 : oai22 port map ( Y=>nx452, A0=>nx9061, A1=>nx9075, B0=>nx9087, B1
      =>nx9089);
   booth_integrtaion_9_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_31, QB=>nx9087, D=>nx3241, CLK=>clk, 
      R=>rst);
   ix9098 : inv01 port map ( Y=>nx9097, A=>weight_9(14));
   ix9102 : aoi22 port map ( Y=>nx9101, A0=>weight_9(15), A1=>nx102, B0=>
      nx106, B1=>nx454);
   ix455 : xnor2 port map ( Y=>nx454, A0=>weight_9(15), A1=>nx438);
   ix439 : nor02ii port map ( Y=>nx438, A0=>weight_9(14), A1=>nx414);
   ix449 : oai32 port map ( Y=>nx448, A0=>nx9109, A1=>nx14402, A2=>nx438, B0
      =>nx9097, B1=>nx14406);
   ix9110 : nor02ii port map ( Y=>nx9109, A0=>nx414, A1=>weight_9(14));
   ix401 : oai32 port map ( Y=>nx400, A0=>nx9113, A1=>nx14404, A2=>nx390, B0
      =>nx9049, B1=>nx14408);
   ix9114 : nor02ii port map ( Y=>nx9113, A0=>nx366, A1=>weight_9(12));
   ix353 : oai32 port map ( Y=>nx352, A0=>nx9117, A1=>nx14404, A2=>nx342, B0
      =>nx9001, B1=>nx14408);
   ix9118 : nor02ii port map ( Y=>nx9117, A0=>nx318, A1=>weight_9(10));
   ix305 : oai32 port map ( Y=>nx304, A0=>nx9121, A1=>nx14404, A2=>nx294, B0
      =>nx8958, B1=>nx14408);
   ix9122 : nor02ii port map ( Y=>nx9121, A0=>nx270, A1=>weight_9(8));
   ix257 : oai32 port map ( Y=>nx256, A0=>nx9125, A1=>nx14404, A2=>nx246, B0
      =>nx8922, B1=>nx14408);
   ix9126 : nor02ii port map ( Y=>nx9125, A0=>nx222, A1=>weight_9(6));
   ix209 : oai32 port map ( Y=>nx208, A0=>nx9129, A1=>nx14404, A2=>nx198, B0
      =>nx8886, B1=>nx14408);
   ix9130 : nor02ii port map ( Y=>nx9129, A0=>nx174, A1=>weight_9(4));
   ix9134 : aoi32 port map ( Y=>nx9133, A0=>nx120, A1=>nx106, A2=>nx8813, B0
      =>weight_9(1), B1=>nx102);
   booth_integrtaion_9_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_9_booth_output_16, QB=>nx8785, D=>nx3381, CLK=>clk, 
      R=>rst);
   booth_integrtaion_9_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_9_15, QB=>nx9139, D=>nx3391, CLK=>clk, R=>rst
   );
   ix985 : xor2 port map ( Y=>label_9(1), A0=>nx9165, A1=>nx9167);
   ix9166 : nand02 port map ( Y=>nx9165, A0=>adderInput_9(0), A1=>
      booth_integration_output_9_0);
   ix9168 : xnor2 port map ( Y=>nx9167, A0=>booth_integration_output_9_1, A1
      =>adderInput_9(1));
   ix983 : xor2 port map ( Y=>label_9(2), A0=>nx9171, A1=>nx9175);
   ix9172 : aoi32 port map ( Y=>nx9171, A0=>adderInput_9(0), A1=>
      booth_integration_output_9_0, A2=>nx842, B0=>adderInput_9(1), B1=>
      booth_integration_output_9_1);
   ix981 : xnor2 port map ( Y=>label_9(3), A0=>nx856, A1=>nx9183);
   ix857 : oai22 port map ( Y=>nx856, A0=>nx9171, A1=>nx9175, B0=>nx9181, B1
      =>nx9161);
   ix9182 : inv01 port map ( Y=>nx9181, A=>adderInput_9(2));
   ix9184 : xnor2 port map ( Y=>nx9183, A0=>booth_integration_output_9_3, A1
      =>adderInput_9(3));
   ix979 : xor2 port map ( Y=>label_9(4), A0=>nx9187, A1=>nx9191);
   ix9188 : aoi22 port map ( Y=>nx9187, A0=>adderInput_9(3), A1=>
      booth_integration_output_9_3, B0=>nx856, B1=>nx858);
   ix977 : xnor2 port map ( Y=>label_9(5), A0=>nx872, A1=>nx9199);
   ix873 : oai22 port map ( Y=>nx872, A0=>nx9187, A1=>nx9191, B0=>nx9197, B1
      =>nx9157);
   ix9198 : inv01 port map ( Y=>nx9197, A=>adderInput_9(4));
   ix9200 : xnor2 port map ( Y=>nx9199, A0=>booth_integration_output_9_5, A1
      =>adderInput_9(5));
   ix975 : xor2 port map ( Y=>label_9(6), A0=>nx9203, A1=>nx9207);
   ix9204 : aoi22 port map ( Y=>nx9203, A0=>adderInput_9(5), A1=>
      booth_integration_output_9_5, B0=>nx872, B1=>nx874);
   ix973 : xnor2 port map ( Y=>label_9(7), A0=>nx888, A1=>nx9215);
   ix889 : oai22 port map ( Y=>nx888, A0=>nx9203, A1=>nx9207, B0=>nx9213, B1
      =>nx9153);
   ix9214 : inv01 port map ( Y=>nx9213, A=>adderInput_9(6));
   ix9216 : xnor2 port map ( Y=>nx9215, A0=>booth_integration_output_9_7, A1
      =>adderInput_9(7));
   ix971 : xor2 port map ( Y=>label_9(8), A0=>nx9219, A1=>nx9223);
   ix9220 : aoi22 port map ( Y=>nx9219, A0=>adderInput_9(7), A1=>
      booth_integration_output_9_7, B0=>nx888, B1=>nx890);
   ix969 : xnor2 port map ( Y=>label_9(9), A0=>nx904, A1=>nx9231);
   ix905 : oai22 port map ( Y=>nx904, A0=>nx9219, A1=>nx9223, B0=>nx9229, B1
      =>nx9149);
   ix9230 : inv01 port map ( Y=>nx9229, A=>adderInput_9(8));
   ix9232 : xnor2 port map ( Y=>nx9231, A0=>booth_integration_output_9_9, A1
      =>adderInput_9(9));
   ix967 : xor2 port map ( Y=>label_9(10), A0=>nx9235, A1=>nx9239);
   ix9236 : aoi22 port map ( Y=>nx9235, A0=>adderInput_9(9), A1=>
      booth_integration_output_9_9, B0=>nx904, B1=>nx906);
   ix965 : xnor2 port map ( Y=>label_9(11), A0=>nx920, A1=>nx9247);
   ix921 : oai22 port map ( Y=>nx920, A0=>nx9235, A1=>nx9239, B0=>nx9245, B1
      =>nx9146);
   ix9246 : inv01 port map ( Y=>nx9245, A=>adderInput_9(10));
   ix9248 : xnor2 port map ( Y=>nx9247, A0=>booth_integration_output_9_11, 
      A1=>adderInput_9(11));
   ix963 : xor2 port map ( Y=>label_9(12), A0=>nx9251, A1=>nx9255);
   ix9252 : aoi22 port map ( Y=>nx9251, A0=>adderInput_9(11), A1=>
      booth_integration_output_9_11, B0=>nx920, B1=>nx922);
   ix961 : xnor2 port map ( Y=>label_9(13), A0=>nx936, A1=>nx9263);
   ix937 : oai22 port map ( Y=>nx936, A0=>nx9251, A1=>nx9255, B0=>nx9261, B1
      =>nx9143);
   ix9262 : inv01 port map ( Y=>nx9261, A=>adderInput_9(12));
   ix9264 : xnor2 port map ( Y=>nx9263, A0=>booth_integration_output_9_13, 
      A1=>adderInput_9(13));
   ix959 : xor2 port map ( Y=>label_9(14), A0=>nx9267, A1=>nx9271);
   ix9268 : aoi22 port map ( Y=>nx9267, A0=>adderInput_9(13), A1=>
      booth_integration_output_9_13, B0=>nx936, B1=>nx938);
   ix957 : xnor2 port map ( Y=>label_9(15), A0=>nx952, A1=>nx9279);
   ix953 : oai22 port map ( Y=>nx952, A0=>nx9267, A1=>nx9271, B0=>nx9277, B1
      =>nx9141);
   ix9278 : inv01 port map ( Y=>nx9277, A=>adderInput_9(14));
   booth_integrtaion_8_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_1, QB=>OPEN, D=>nx4061, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_2, QB=>nx9833, D=>nx4051, CLK=>clk, R=>rst
   );
   booth_integrtaion_8_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_3, QB=>OPEN, D=>nx4041, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_4, QB=>nx9831, D=>nx4031, CLK=>clk, R=>rst
   );
   booth_integrtaion_8_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_5, QB=>OPEN, D=>nx4021, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_6, QB=>nx9829, D=>nx4011, CLK=>clk, R=>rst
   );
   booth_integrtaion_8_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_7, QB=>OPEN, D=>nx4001, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_8, QB=>nx9825, D=>nx3991, CLK=>clk, R=>rst
   );
   booth_integrtaion_8_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_9, QB=>OPEN, D=>nx3981, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_10, QB=>nx9821, D=>nx3971, CLK=>clk, R=>rst
   );
   booth_integrtaion_8_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_11, QB=>OPEN, D=>nx3961, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_12, QB=>nx9817, D=>nx3951, CLK=>clk, R=>rst
   );
   booth_integrtaion_8_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_13, QB=>OPEN, D=>nx3941, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_14, QB=>nx9813, D=>nx3931, CLK=>clk, R=>rst
   );
   ix9362 : aoi22 port map ( Y=>nx9361, A0=>neuron(15), A1=>nx14196, B0=>
      nx1628, B1=>nx1634);
   booth_integrtaion_8_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_reg_output_0, QB=>OPEN, D=>nx3571, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_0, QB=>OPEN, D=>nx3557, CLK=>clk, 
      S=>nx14146);
   booth_integrtaion_8_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_reg_output_9, QB=>OPEN, D=>nx3751, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_9, QB=>OPEN, D=>nx3741, CLK=>clk, 
      R=>nx14146);
   booth_integrtaion_8_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_8, QB=>OPEN, D=>nx3731, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_8, QB=>OPEN, D=>nx3721, CLK=>clk, 
      R=>nx14146);
   booth_integrtaion_8_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_7, QB=>OPEN, D=>nx3711, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_7, QB=>OPEN, D=>nx3701, CLK=>clk, 
      R=>nx14146);
   booth_integrtaion_8_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_6, QB=>OPEN, D=>nx3691, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_6, QB=>OPEN, D=>nx3681, CLK=>clk, 
      R=>nx14146);
   booth_integrtaion_8_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_5, QB=>OPEN, D=>nx3671, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_5, QB=>OPEN, D=>nx3661, CLK=>clk, 
      R=>nx14146);
   booth_integrtaion_8_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_4, QB=>OPEN, D=>nx3651, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_4, QB=>OPEN, D=>nx3641, CLK=>clk, 
      R=>nx14146);
   booth_integrtaion_8_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_3, QB=>OPEN, D=>nx3631, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_3, QB=>OPEN, D=>nx3621, CLK=>clk, 
      R=>nx14144);
   booth_integrtaion_8_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_2, QB=>OPEN, D=>nx3611, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_2, QB=>OPEN, D=>nx3601, CLK=>clk, 
      R=>nx14144);
   booth_integrtaion_8_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_output_1, QB=>OPEN, D=>nx3591, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_8_shift_Reg_count_1, QB=>OPEN, D=>nx3581, CLK=>clk, 
      R=>nx14144);
   ix3552 : nand02 port map ( Y=>nx3551, A0=>nx14616, A1=>nx14182);
   booth_integrtaion_8_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx9423, D=>nx3551, CLK=>clk, S=>nx14144);
   ix1629 : nand02 port map ( Y=>nx1628, A0=>nx9447, A1=>nx9461);
   ix9448 : oai21 port map ( Y=>nx9447, A0=>nx1092, A1=>nx1088, B0=>
      weight_8(0));
   ix3762 : oai21 port map ( Y=>nx3761, A0=>nx9453, A1=>nx14410, B0=>nx9455
   );
   booth_integrtaion_8_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9453, D=>nx3761, CLK=>clk, R=>rst);
   booth_integrtaion_8_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_0, QB=>nx9283, D=>nx4071, CLK=>clk, R=>rst
   );
   ix9467 : xnor2 port map ( Y=>nx9466, A0=>nx1098, A1=>nx2831);
   ix3902 : oai21 port map ( Y=>nx3901, A0=>nx9475, A1=>nx14410, B0=>nx9477
   );
   booth_integrtaion_8_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_17, QB=>nx9475, D=>nx3901, CLK=>clk, 
      R=>rst);
   ix9478 : nand03 port map ( Y=>nx9477, A0=>nx14418, A1=>nx1606, A2=>
      nx14674);
   ix1607 : xnor2 port map ( Y=>nx1606, A0=>nx9480, A1=>nx2833);
   ix9482 : aoi22 port map ( Y=>nx9480, A0=>
      booth_integrtaion_8_booth_output_17, A1=>nx1122, B0=>nx1098, B1=>
      nx2831);
   ix1107 : nand02 port map ( Y=>nx1106, A0=>weight_8(1), A1=>weight_8(0));
   ix9488 : or02 port map ( Y=>nx9487, A0=>weight_8(0), A1=>weight_8(1));
   ix3892 : oai21 port map ( Y=>nx3891, A0=>nx9492, A1=>nx14410, B0=>nx9495
   );
   booth_integrtaion_8_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9492, D=>nx3891, CLK=>clk, R=>rst);
   ix9496 : nand03 port map ( Y=>nx9495, A0=>nx14418, A1=>nx1594, A2=>
      nx14674);
   ix1595 : xnor2 port map ( Y=>nx1594, A0=>nx1150, A1=>nx9507);
   ix1151 : oai22 port map ( Y=>nx1150, A0=>nx9480, A1=>nx9499, B0=>nx9492, 
      B1=>nx14422);
   ix9502 : aoi32 port map ( Y=>nx9501, A0=>nx1132, A1=>nx1092, A2=>nx9504, 
      B0=>weight_8(2), B1=>nx1088);
   ix1133 : oai21 port map ( Y=>nx1132, A0=>weight_8(0), A1=>weight_8(1), B0
      =>weight_8(2));
   ix9508 : xnor2 port map ( Y=>nx9507, A0=>
      booth_integrtaion_8_booth_output_19, A1=>nx1170);
   booth_integrtaion_8_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_19, QB=>OPEN, D=>nx3881, CLK=>clk, R
      =>rst);
   ix9514 : xnor2 port map ( Y=>nx9513, A0=>nx9515, A1=>nx9532);
   ix9516 : aoi22 port map ( Y=>nx9515, A0=>
      booth_integrtaion_8_booth_output_19, A1=>nx1170, B0=>nx1150, B1=>
      nx2835);
   ix1171 : oai32 port map ( Y=>nx1170, A0=>nx9519, A1=>nx14424, A2=>nx1160, 
      B0=>nx9527, B1=>nx14428);
   ix9520 : nor02ii port map ( Y=>nx9519, A0=>nx1136, A1=>weight_8(3));
   ix1137 : nor03_2x port map ( Y=>nx1136, A0=>weight_8(2), A1=>weight_8(0), 
      A2=>weight_8(1));
   ix1161 : nor04 port map ( Y=>nx1160, A0=>weight_8(3), A1=>weight_8(2), A2
      =>weight_8(0), A3=>weight_8(1));
   ix9528 : inv01 port map ( Y=>nx9527, A=>weight_8(3));
   ix3872 : oai21 port map ( Y=>nx3871, A0=>nx9537, A1=>nx14410, B0=>nx9539
   );
   booth_integrtaion_8_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9537, D=>nx3871, CLK=>clk, R=>rst);
   ix9540 : nand03 port map ( Y=>nx9539, A0=>nx14418, A1=>nx1570, A2=>
      nx14674);
   ix1571 : xnor2 port map ( Y=>nx1570, A0=>nx1198, A1=>nx9553);
   ix1199 : oai22 port map ( Y=>nx1198, A0=>nx9515, A1=>nx9532, B0=>nx9537, 
      B1=>nx9544);
   ix9552 : inv01 port map ( Y=>nx9551, A=>weight_8(4));
   ix9554 : xnor2 port map ( Y=>nx9553, A0=>
      booth_integrtaion_8_booth_output_21, A1=>nx1218);
   booth_integrtaion_8_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_21, QB=>OPEN, D=>nx3861, CLK=>clk, R
      =>rst);
   ix9559 : xnor2 port map ( Y=>nx9558, A0=>nx9561, A1=>nx9573);
   ix9562 : aoi22 port map ( Y=>nx9561, A0=>
      booth_integrtaion_8_booth_output_21, A1=>nx1218, B0=>nx1198, B1=>
      nx2839);
   ix1219 : oai32 port map ( Y=>nx1218, A0=>nx9565, A1=>nx14424, A2=>nx1208, 
      B0=>nx9569, B1=>nx14428);
   ix9566 : nor02ii port map ( Y=>nx9565, A0=>nx1184, A1=>weight_8(5));
   ix1185 : nor02ii port map ( Y=>nx1184, A0=>weight_8(4), A1=>nx1160);
   ix1209 : nor02ii port map ( Y=>nx1208, A0=>weight_8(5), A1=>nx1184);
   ix9570 : inv01 port map ( Y=>nx9569, A=>weight_8(5));
   ix3852 : oai21 port map ( Y=>nx3851, A0=>nx9579, A1=>nx14410, B0=>nx9581
   );
   booth_integrtaion_8_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9579, D=>nx3851, CLK=>clk, R=>rst);
   ix9582 : nand03 port map ( Y=>nx9581, A0=>nx14418, A1=>nx1546, A2=>
      nx14412);
   ix1547 : xnor2 port map ( Y=>nx1546, A0=>nx1246, A1=>nx9595);
   ix1247 : oai22 port map ( Y=>nx1246, A0=>nx9561, A1=>nx9573, B0=>nx9579, 
      B1=>nx9585);
   ix9594 : inv01 port map ( Y=>nx9593, A=>weight_8(6));
   ix9596 : xnor2 port map ( Y=>nx9595, A0=>
      booth_integrtaion_8_booth_output_23, A1=>nx1266);
   booth_integrtaion_8_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_23, QB=>OPEN, D=>nx3841, CLK=>clk, R
      =>rst);
   ix9604 : xnor2 port map ( Y=>nx9603, A0=>nx9605, A1=>nx9618);
   ix9606 : aoi22 port map ( Y=>nx9605, A0=>
      booth_integrtaion_8_booth_output_23, A1=>nx1266, B0=>nx1246, B1=>
      nx2843);
   ix1267 : oai32 port map ( Y=>nx1266, A0=>nx9609, A1=>nx14424, A2=>nx1256, 
      B0=>nx9615, B1=>nx14428);
   ix9610 : nor02ii port map ( Y=>nx9609, A0=>nx1232, A1=>weight_8(7));
   ix1233 : nor02ii port map ( Y=>nx1232, A0=>weight_8(6), A1=>nx1208);
   ix1257 : nor02ii port map ( Y=>nx1256, A0=>weight_8(7), A1=>nx1232);
   ix9616 : inv01 port map ( Y=>nx9615, A=>weight_8(7));
   ix3832 : oai21 port map ( Y=>nx3831, A0=>nx9623, A1=>nx14412, B0=>nx9625
   );
   booth_integrtaion_8_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9623, D=>nx3831, CLK=>clk, R=>rst);
   ix9626 : nand03 port map ( Y=>nx9625, A0=>nx14418, A1=>nx1522, A2=>
      nx14412);
   ix1523 : xnor2 port map ( Y=>nx1522, A0=>nx1294, A1=>nx9639);
   ix1295 : oai22 port map ( Y=>nx1294, A0=>nx9605, A1=>nx9618, B0=>nx9623, 
      B1=>nx9629);
   ix9638 : inv01 port map ( Y=>nx9637, A=>weight_8(8));
   ix9640 : xnor2 port map ( Y=>nx9639, A0=>
      booth_integrtaion_8_booth_output_25, A1=>nx1314);
   booth_integrtaion_8_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_25, QB=>OPEN, D=>nx3821, CLK=>clk, R
      =>rst);
   ix9646 : xnor2 port map ( Y=>nx9645, A0=>nx9647, A1=>nx9659);
   ix9648 : aoi22 port map ( Y=>nx9647, A0=>
      booth_integrtaion_8_booth_output_25, A1=>nx1314, B0=>nx1294, B1=>
      nx2847);
   ix1315 : oai32 port map ( Y=>nx1314, A0=>nx9651, A1=>nx14424, A2=>nx1304, 
      B0=>nx9655, B1=>nx14428);
   ix9652 : nor02ii port map ( Y=>nx9651, A0=>nx1280, A1=>weight_8(9));
   ix1281 : nor02ii port map ( Y=>nx1280, A0=>weight_8(8), A1=>nx1256);
   ix1305 : nor02ii port map ( Y=>nx1304, A0=>weight_8(9), A1=>nx1280);
   ix9656 : inv01 port map ( Y=>nx9655, A=>weight_8(9));
   ix3812 : oai21 port map ( Y=>nx3811, A0=>nx9664, A1=>nx14412, B0=>nx9666
   );
   booth_integrtaion_8_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9664, D=>nx3811, CLK=>clk, R=>rst);
   ix9667 : nand03 port map ( Y=>nx9666, A0=>nx14418, A1=>nx1498, A2=>
      nx14412);
   ix1499 : xnor2 port map ( Y=>nx1498, A0=>nx1342, A1=>nx9681);
   ix1343 : oai22 port map ( Y=>nx1342, A0=>nx9647, A1=>nx9659, B0=>nx9664, 
      B1=>nx9671);
   ix9680 : inv01 port map ( Y=>nx9679, A=>weight_8(10));
   ix9682 : xnor2 port map ( Y=>nx9681, A0=>
      booth_integrtaion_8_booth_output_27, A1=>nx1362);
   booth_integrtaion_8_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_27, QB=>OPEN, D=>nx3801, CLK=>clk, R
      =>rst);
   ix9689 : xnor2 port map ( Y=>nx9688, A0=>nx9690, A1=>nx9702);
   ix9691 : aoi22 port map ( Y=>nx9690, A0=>
      booth_integrtaion_8_booth_output_27, A1=>nx1362, B0=>nx1342, B1=>
      nx2851);
   ix1363 : oai32 port map ( Y=>nx1362, A0=>nx9693, A1=>nx14424, A2=>nx1352, 
      B0=>nx9699, B1=>nx14428);
   ix9694 : nor02ii port map ( Y=>nx9693, A0=>nx1328, A1=>weight_8(11));
   ix1329 : nor02ii port map ( Y=>nx1328, A0=>weight_8(10), A1=>nx1304);
   ix1353 : nor02ii port map ( Y=>nx1352, A0=>weight_8(11), A1=>nx1328);
   ix9700 : inv01 port map ( Y=>nx9699, A=>weight_8(11));
   ix3792 : oai21 port map ( Y=>nx3791, A0=>nx9707, A1=>nx14412, B0=>nx9709
   );
   booth_integrtaion_8_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx9707, D=>nx3791, CLK=>clk, R=>rst);
   ix9710 : nand03 port map ( Y=>nx9709, A0=>nx14682, A1=>nx1474, A2=>
      nx14412);
   ix1475 : xnor2 port map ( Y=>nx1474, A0=>nx1390, A1=>nx9723);
   ix1391 : oai22 port map ( Y=>nx1390, A0=>nx9690, A1=>nx9702, B0=>nx9707, 
      B1=>nx9713);
   ix9722 : inv01 port map ( Y=>nx9721, A=>weight_8(12));
   ix9724 : xnor2 port map ( Y=>nx9723, A0=>
      booth_integrtaion_8_booth_output_29, A1=>nx1410);
   booth_integrtaion_8_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_29, QB=>OPEN, D=>nx3781, CLK=>clk, R
      =>rst);
   ix9732 : xnor2 port map ( Y=>nx9731, A0=>nx9733, A1=>nx9747);
   ix9734 : aoi22 port map ( Y=>nx9733, A0=>
      booth_integrtaion_8_booth_output_29, A1=>nx1410, B0=>nx1390, B1=>
      nx2855);
   ix1411 : oai32 port map ( Y=>nx1410, A0=>nx9737, A1=>nx14424, A2=>nx1400, 
      B0=>nx9743, B1=>nx14428);
   ix9738 : nor02ii port map ( Y=>nx9737, A0=>nx1376, A1=>weight_8(13));
   ix1377 : nor02ii port map ( Y=>nx1376, A0=>weight_8(12), A1=>nx1352);
   ix1401 : nor02ii port map ( Y=>nx1400, A0=>weight_8(13), A1=>nx1376);
   ix9744 : inv01 port map ( Y=>nx9743, A=>weight_8(13));
   ix9756 : xnor2 port map ( Y=>nx9755, A0=>nx1438, A1=>nx1448);
   ix1439 : oai22 port map ( Y=>nx1438, A0=>nx9733, A1=>nx9747, B0=>nx9759, 
      B1=>nx9761);
   booth_integrtaion_8_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_31, QB=>nx9759, D=>nx3771, CLK=>clk, 
      R=>rst);
   ix9770 : inv01 port map ( Y=>nx9769, A=>weight_8(14));
   ix9774 : aoi22 port map ( Y=>nx9773, A0=>weight_8(15), A1=>nx1088, B0=>
      nx1092, B1=>nx1440);
   ix1441 : xnor2 port map ( Y=>nx1440, A0=>weight_8(15), A1=>nx1424);
   ix1425 : nor02ii port map ( Y=>nx1424, A0=>weight_8(14), A1=>nx1400);
   ix1435 : oai32 port map ( Y=>nx1434, A0=>nx9781, A1=>nx14424, A2=>nx1424, 
      B0=>nx9769, B1=>nx14428);
   ix9782 : nor02ii port map ( Y=>nx9781, A0=>nx1400, A1=>weight_8(14));
   ix1387 : oai32 port map ( Y=>nx1386, A0=>nx9785, A1=>nx14426, A2=>nx1376, 
      B0=>nx9721, B1=>nx14430);
   ix9786 : nor02ii port map ( Y=>nx9785, A0=>nx1352, A1=>weight_8(12));
   ix1339 : oai32 port map ( Y=>nx1338, A0=>nx9789, A1=>nx14426, A2=>nx1328, 
      B0=>nx9679, B1=>nx14430);
   ix9790 : nor02ii port map ( Y=>nx9789, A0=>nx1304, A1=>weight_8(10));
   ix1291 : oai32 port map ( Y=>nx1290, A0=>nx9793, A1=>nx14426, A2=>nx1280, 
      B0=>nx9637, B1=>nx14430);
   ix9794 : nor02ii port map ( Y=>nx9793, A0=>nx1256, A1=>weight_8(8));
   ix1243 : oai32 port map ( Y=>nx1242, A0=>nx9797, A1=>nx14426, A2=>nx1232, 
      B0=>nx9593, B1=>nx14430);
   ix9798 : nor02ii port map ( Y=>nx9797, A0=>nx1208, A1=>weight_8(6));
   ix1195 : oai32 port map ( Y=>nx1194, A0=>nx9801, A1=>nx14426, A2=>nx1184, 
      B0=>nx9551, B1=>nx14430);
   ix9802 : nor02ii port map ( Y=>nx9801, A0=>nx1160, A1=>weight_8(4));
   ix9806 : aoi32 port map ( Y=>nx9805, A0=>nx1106, A1=>nx1092, A2=>nx9487, 
      B0=>weight_8(1), B1=>nx1088);
   booth_integrtaion_8_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_8_booth_output_16, QB=>nx9461, D=>nx3911, CLK=>clk, 
      R=>rst);
   booth_integrtaion_8_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_8_15, QB=>nx9811, D=>nx3921, CLK=>clk, R=>rst
   );
   ix1971 : xor2 port map ( Y=>label_8(1), A0=>nx9837, A1=>nx9839);
   ix9838 : nand02 port map ( Y=>nx9837, A0=>adderInput_8(0), A1=>
      booth_integration_output_8_0);
   ix9840 : xnor2 port map ( Y=>nx9839, A0=>booth_integration_output_8_1, A1
      =>adderInput_8(1));
   ix1969 : xor2 port map ( Y=>label_8(2), A0=>nx9843, A1=>nx9847);
   ix9844 : aoi32 port map ( Y=>nx9843, A0=>adderInput_8(0), A1=>
      booth_integration_output_8_0, A2=>nx1828, B0=>adderInput_8(1), B1=>
      booth_integration_output_8_1);
   ix1967 : xnor2 port map ( Y=>label_8(3), A0=>nx1842, A1=>nx9855);
   ix1843 : oai22 port map ( Y=>nx1842, A0=>nx9843, A1=>nx9847, B0=>nx9853, 
      B1=>nx9833);
   ix9854 : inv01 port map ( Y=>nx9853, A=>adderInput_8(2));
   ix9856 : xnor2 port map ( Y=>nx9855, A0=>booth_integration_output_8_3, A1
      =>adderInput_8(3));
   ix1965 : xor2 port map ( Y=>label_8(4), A0=>nx9859, A1=>nx9863);
   ix9860 : aoi22 port map ( Y=>nx9859, A0=>adderInput_8(3), A1=>
      booth_integration_output_8_3, B0=>nx1842, B1=>nx1844);
   ix1963 : xnor2 port map ( Y=>label_8(5), A0=>nx1858, A1=>nx9870);
   ix1859 : oai22 port map ( Y=>nx1858, A0=>nx9859, A1=>nx9863, B0=>nx9868, 
      B1=>nx9831);
   ix9869 : inv01 port map ( Y=>nx9868, A=>adderInput_8(4));
   ix9872 : xnor2 port map ( Y=>nx9870, A0=>booth_integration_output_8_5, A1
      =>adderInput_8(5));
   ix1961 : xor2 port map ( Y=>label_8(6), A0=>nx9874, A1=>nx9877);
   ix9875 : aoi22 port map ( Y=>nx9874, A0=>adderInput_8(5), A1=>
      booth_integration_output_8_5, B0=>nx1858, B1=>nx1860);
   ix1959 : xnor2 port map ( Y=>label_8(7), A0=>nx1874, A1=>nx9883);
   ix1875 : oai22 port map ( Y=>nx1874, A0=>nx9874, A1=>nx9877, B0=>nx9881, 
      B1=>nx9829);
   ix9882 : inv01 port map ( Y=>nx9881, A=>adderInput_8(6));
   ix9884 : xnor2 port map ( Y=>nx9883, A0=>booth_integration_output_8_7, A1
      =>adderInput_8(7));
   ix1957 : xor2 port map ( Y=>label_8(8), A0=>nx9886, A1=>nx9889);
   ix9887 : aoi22 port map ( Y=>nx9886, A0=>adderInput_8(7), A1=>
      booth_integration_output_8_7, B0=>nx1874, B1=>nx1876);
   ix1955 : xnor2 port map ( Y=>label_8(9), A0=>nx1890, A1=>nx9895);
   ix1891 : oai22 port map ( Y=>nx1890, A0=>nx9886, A1=>nx9889, B0=>nx9893, 
      B1=>nx9825);
   ix9894 : inv01 port map ( Y=>nx9893, A=>adderInput_8(8));
   ix9896 : xnor2 port map ( Y=>nx9895, A0=>booth_integration_output_8_9, A1
      =>adderInput_8(9));
   ix1953 : xor2 port map ( Y=>label_8(10), A0=>nx9898, A1=>nx9901);
   ix9899 : aoi22 port map ( Y=>nx9898, A0=>adderInput_8(9), A1=>
      booth_integration_output_8_9, B0=>nx1890, B1=>nx1892);
   ix1951 : xnor2 port map ( Y=>label_8(11), A0=>nx1906, A1=>nx9907);
   ix1907 : oai22 port map ( Y=>nx1906, A0=>nx9898, A1=>nx9901, B0=>nx9905, 
      B1=>nx9821);
   ix9906 : inv01 port map ( Y=>nx9905, A=>adderInput_8(10));
   ix9908 : xnor2 port map ( Y=>nx9907, A0=>booth_integration_output_8_11, 
      A1=>adderInput_8(11));
   ix1949 : xor2 port map ( Y=>label_8(12), A0=>nx9910, A1=>nx9913);
   ix9911 : aoi22 port map ( Y=>nx9910, A0=>adderInput_8(11), A1=>
      booth_integration_output_8_11, B0=>nx1906, B1=>nx1908);
   ix1947 : xnor2 port map ( Y=>label_8(13), A0=>nx1922, A1=>nx9919);
   ix1923 : oai22 port map ( Y=>nx1922, A0=>nx9910, A1=>nx9913, B0=>nx9917, 
      B1=>nx9817);
   ix9918 : inv01 port map ( Y=>nx9917, A=>adderInput_8(12));
   ix9920 : xnor2 port map ( Y=>nx9919, A0=>booth_integration_output_8_13, 
      A1=>adderInput_8(13));
   ix1945 : xor2 port map ( Y=>label_8(14), A0=>nx9922, A1=>nx9925);
   ix9923 : aoi22 port map ( Y=>nx9922, A0=>adderInput_8(13), A1=>
      booth_integration_output_8_13, B0=>nx1922, B1=>nx1924);
   ix1943 : xnor2 port map ( Y=>label_8(15), A0=>nx1938, A1=>nx9931);
   ix1939 : oai22 port map ( Y=>nx1938, A0=>nx9922, A1=>nx9925, B0=>nx9929, 
      B1=>nx9813);
   ix9930 : inv01 port map ( Y=>nx9929, A=>adderInput_8(14));
   booth_integrtaion_7_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_1, QB=>OPEN, D=>nx4591, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_2, QB=>nx10365, D=>nx4581, CLK=>clk, R=>rst
   );
   booth_integrtaion_7_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_3, QB=>OPEN, D=>nx4571, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_4, QB=>nx10363, D=>nx4561, CLK=>clk, R=>rst
   );
   booth_integrtaion_7_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_5, QB=>OPEN, D=>nx4551, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_6, QB=>nx10361, D=>nx4541, CLK=>clk, R=>rst
   );
   booth_integrtaion_7_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_7, QB=>OPEN, D=>nx4531, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_8, QB=>nx10359, D=>nx4521, CLK=>clk, R=>rst
   );
   booth_integrtaion_7_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_9, QB=>OPEN, D=>nx4511, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_10, QB=>nx10357, D=>nx4501, CLK=>clk, R=>
      rst);
   booth_integrtaion_7_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_11, QB=>OPEN, D=>nx4491, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_12, QB=>nx10355, D=>nx4481, CLK=>clk, R=>
      rst);
   booth_integrtaion_7_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_13, QB=>OPEN, D=>nx4471, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_14, QB=>nx10353, D=>nx4461, CLK=>clk, R=>
      rst);
   ix9983 : aoi22 port map ( Y=>nx9982, A0=>neuron(15), A1=>nx14218, B0=>
      nx2614, B1=>nx2620);
   booth_integrtaion_7_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_reg_output_0, QB=>OPEN, D=>nx4101, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_0, QB=>OPEN, D=>nx4087, CLK=>clk, 
      S=>nx14150);
   booth_integrtaion_7_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_reg_output_9, QB=>OPEN, D=>nx4281, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_9, QB=>OPEN, D=>nx4271, CLK=>clk, 
      R=>nx14150);
   booth_integrtaion_7_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_8, QB=>OPEN, D=>nx4261, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_8, QB=>OPEN, D=>nx4251, CLK=>clk, 
      R=>nx14150);
   booth_integrtaion_7_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_7, QB=>OPEN, D=>nx4241, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_7, QB=>OPEN, D=>nx4231, CLK=>clk, 
      R=>nx14150);
   booth_integrtaion_7_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_6, QB=>OPEN, D=>nx4221, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_6, QB=>OPEN, D=>nx4211, CLK=>clk, 
      R=>nx14148);
   booth_integrtaion_7_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_5, QB=>OPEN, D=>nx4201, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_5, QB=>OPEN, D=>nx4191, CLK=>clk, 
      R=>nx14148);
   booth_integrtaion_7_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_4, QB=>OPEN, D=>nx4181, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_4, QB=>OPEN, D=>nx4171, CLK=>clk, 
      R=>nx14148);
   booth_integrtaion_7_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_3, QB=>OPEN, D=>nx4161, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_3, QB=>OPEN, D=>nx4151, CLK=>clk, 
      R=>nx14148);
   booth_integrtaion_7_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_2, QB=>OPEN, D=>nx4141, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_2, QB=>OPEN, D=>nx4131, CLK=>clk, 
      R=>nx14148);
   booth_integrtaion_7_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_output_1, QB=>OPEN, D=>nx4121, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_7_shift_Reg_count_1, QB=>OPEN, D=>nx4111, CLK=>clk, 
      R=>nx14148);
   ix4082 : nand02 port map ( Y=>nx4081, A0=>nx14620, A1=>nx14204);
   booth_integrtaion_7_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx10029, D=>nx4081, CLK=>clk, S=>nx14148);
   ix2615 : nand02 port map ( Y=>nx2614, A0=>nx10050, A1=>nx10061);
   ix10051 : oai21 port map ( Y=>nx10050, A0=>nx2078, A1=>nx2074, B0=>
      weight_7(0));
   ix4292 : oai21 port map ( Y=>nx4291, A0=>nx10055, A1=>nx14432, B0=>
      nx10057);
   booth_integrtaion_7_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10055, D=>nx4291, CLK=>clk, R=>rst);
   booth_integrtaion_7_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_0, QB=>nx9934, D=>nx4601, CLK=>clk, R=>rst
   );
   ix10066 : xnor2 port map ( Y=>nx10065, A0=>nx2084, A1=>nx2861);
   ix4432 : oai21 port map ( Y=>nx4431, A0=>nx10071, A1=>nx14432, B0=>
      nx10073);
   booth_integrtaion_7_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_17, QB=>nx10071, D=>nx4431, CLK=>clk, 
      R=>rst);
   ix10074 : nand03 port map ( Y=>nx10073, A0=>nx14440, A1=>nx2592, A2=>
      nx14690);
   ix2593 : xnor2 port map ( Y=>nx2592, A0=>nx10076, A1=>nx2863);
   ix10077 : aoi22 port map ( Y=>nx10076, A0=>
      booth_integrtaion_7_booth_output_17, A1=>nx2108, B0=>nx2084, B1=>
      nx2861);
   ix2093 : nand02 port map ( Y=>nx2092, A0=>weight_7(1), A1=>weight_7(0));
   ix10081 : or02 port map ( Y=>nx10080, A0=>weight_7(0), A1=>weight_7(1));
   ix4422 : oai21 port map ( Y=>nx4421, A0=>nx10085, A1=>nx14432, B0=>
      nx10087);
   booth_integrtaion_7_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10085, D=>nx4421, CLK=>clk, R=>rst);
   ix10088 : nand03 port map ( Y=>nx10087, A0=>nx14440, A1=>nx2580, A2=>
      nx14690);
   ix2581 : xnor2 port map ( Y=>nx2580, A0=>nx2136, A1=>nx10098);
   ix2137 : oai22 port map ( Y=>nx2136, A0=>nx10076, A1=>nx10091, B0=>
      nx10085, B1=>nx14444);
   ix10094 : aoi32 port map ( Y=>nx10093, A0=>nx2118, A1=>nx2078, A2=>
      nx10096, B0=>weight_7(2), B1=>nx2074);
   ix2119 : oai21 port map ( Y=>nx2118, A0=>weight_7(0), A1=>weight_7(1), B0
      =>weight_7(2));
   ix10099 : xnor2 port map ( Y=>nx10098, A0=>
      booth_integrtaion_7_booth_output_19, A1=>nx2156);
   booth_integrtaion_7_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_19, QB=>OPEN, D=>nx4411, CLK=>clk, R
      =>rst);
   ix10104 : xnor2 port map ( Y=>nx10103, A0=>nx10105, A1=>nx10119);
   ix10106 : aoi22 port map ( Y=>nx10105, A0=>
      booth_integrtaion_7_booth_output_19, A1=>nx2156, B0=>nx2136, B1=>
      nx2865);
   ix2157 : oai32 port map ( Y=>nx2156, A0=>nx10108, A1=>nx14446, A2=>nx2146, 
      B0=>nx10114, B1=>nx14450);
   ix10109 : nor02ii port map ( Y=>nx10108, A0=>nx2122, A1=>weight_7(3));
   ix2123 : nor03_2x port map ( Y=>nx2122, A0=>weight_7(2), A1=>weight_7(0), 
      A2=>weight_7(1));
   ix2147 : nor04 port map ( Y=>nx2146, A0=>weight_7(3), A1=>weight_7(2), A2
      =>weight_7(0), A3=>weight_7(1));
   ix10115 : inv01 port map ( Y=>nx10114, A=>weight_7(3));
   ix4402 : oai21 port map ( Y=>nx4401, A0=>nx10123, A1=>nx14432, B0=>
      nx10125);
   booth_integrtaion_7_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10123, D=>nx4401, CLK=>clk, R=>rst);
   ix10126 : nand03 port map ( Y=>nx10125, A0=>nx14440, A1=>nx2556, A2=>
      nx14690);
   ix2557 : xnor2 port map ( Y=>nx2556, A0=>nx2184, A1=>nx10138);
   ix2185 : oai22 port map ( Y=>nx2184, A0=>nx10105, A1=>nx10119, B0=>
      nx10123, B1=>nx10129);
   ix10137 : inv01 port map ( Y=>nx10136, A=>weight_7(4));
   ix10139 : xnor2 port map ( Y=>nx10138, A0=>
      booth_integrtaion_7_booth_output_21, A1=>nx2204);
   booth_integrtaion_7_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_21, QB=>OPEN, D=>nx4391, CLK=>clk, R
      =>rst);
   ix10144 : xnor2 port map ( Y=>nx10143, A0=>nx10145, A1=>nx10155);
   ix10146 : aoi22 port map ( Y=>nx10145, A0=>
      booth_integrtaion_7_booth_output_21, A1=>nx2204, B0=>nx2184, B1=>
      nx2869);
   ix2205 : oai32 port map ( Y=>nx2204, A0=>nx10148, A1=>nx14446, A2=>nx2194, 
      B0=>nx10152, B1=>nx14450);
   ix10149 : nor02ii port map ( Y=>nx10148, A0=>nx2170, A1=>weight_7(5));
   ix2171 : nor02ii port map ( Y=>nx2170, A0=>weight_7(4), A1=>nx2146);
   ix2195 : nor02ii port map ( Y=>nx2194, A0=>weight_7(5), A1=>nx2170);
   ix10153 : inv01 port map ( Y=>nx10152, A=>weight_7(5));
   ix4382 : oai21 port map ( Y=>nx4381, A0=>nx10159, A1=>nx14432, B0=>
      nx10161);
   booth_integrtaion_7_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10159, D=>nx4381, CLK=>clk, R=>rst);
   ix10162 : nand03 port map ( Y=>nx10161, A0=>nx14440, A1=>nx2532, A2=>
      nx14434);
   ix2533 : xnor2 port map ( Y=>nx2532, A0=>nx2232, A1=>nx10174);
   ix2233 : oai22 port map ( Y=>nx2232, A0=>nx10145, A1=>nx10155, B0=>
      nx10159, B1=>nx10165);
   ix10173 : inv01 port map ( Y=>nx10172, A=>weight_7(6));
   ix10175 : xnor2 port map ( Y=>nx10174, A0=>
      booth_integrtaion_7_booth_output_23, A1=>nx2252);
   booth_integrtaion_7_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_23, QB=>OPEN, D=>nx4371, CLK=>clk, R
      =>rst);
   ix10180 : xnor2 port map ( Y=>nx10179, A0=>nx10181, A1=>nx10191);
   ix10182 : aoi22 port map ( Y=>nx10181, A0=>
      booth_integrtaion_7_booth_output_23, A1=>nx2252, B0=>nx2232, B1=>
      nx2873);
   ix2253 : oai32 port map ( Y=>nx2252, A0=>nx10184, A1=>nx14446, A2=>nx2242, 
      B0=>nx10188, B1=>nx14450);
   ix10185 : nor02ii port map ( Y=>nx10184, A0=>nx2218, A1=>weight_7(7));
   ix2219 : nor02ii port map ( Y=>nx2218, A0=>weight_7(6), A1=>nx2194);
   ix2243 : nor02ii port map ( Y=>nx2242, A0=>weight_7(7), A1=>nx2218);
   ix10189 : inv01 port map ( Y=>nx10188, A=>weight_7(7));
   ix4362 : oai21 port map ( Y=>nx4361, A0=>nx10195, A1=>nx14434, B0=>
      nx10197);
   booth_integrtaion_7_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10195, D=>nx4361, CLK=>clk, R=>rst);
   ix10198 : nand03 port map ( Y=>nx10197, A0=>nx14440, A1=>nx2508, A2=>
      nx14434);
   ix2509 : xnor2 port map ( Y=>nx2508, A0=>nx2280, A1=>nx10210);
   ix2281 : oai22 port map ( Y=>nx2280, A0=>nx10181, A1=>nx10191, B0=>
      nx10195, B1=>nx10201);
   ix10209 : inv01 port map ( Y=>nx10208, A=>weight_7(8));
   ix10211 : xnor2 port map ( Y=>nx10210, A0=>
      booth_integrtaion_7_booth_output_25, A1=>nx2300);
   booth_integrtaion_7_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_25, QB=>OPEN, D=>nx4351, CLK=>clk, R
      =>rst);
   ix10216 : xnor2 port map ( Y=>nx10215, A0=>nx10217, A1=>nx10227);
   ix10218 : aoi22 port map ( Y=>nx10217, A0=>
      booth_integrtaion_7_booth_output_25, A1=>nx2300, B0=>nx2280, B1=>
      nx2877);
   ix2301 : oai32 port map ( Y=>nx2300, A0=>nx10220, A1=>nx14446, A2=>nx2290, 
      B0=>nx10224, B1=>nx14450);
   ix10221 : nor02ii port map ( Y=>nx10220, A0=>nx2266, A1=>weight_7(9));
   ix2267 : nor02ii port map ( Y=>nx2266, A0=>weight_7(8), A1=>nx2242);
   ix2291 : nor02ii port map ( Y=>nx2290, A0=>weight_7(9), A1=>nx2266);
   ix10225 : inv01 port map ( Y=>nx10224, A=>weight_7(9));
   ix4342 : oai21 port map ( Y=>nx4341, A0=>nx10231, A1=>nx14434, B0=>
      nx10233);
   booth_integrtaion_7_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10231, D=>nx4341, CLK=>clk, R=>rst);
   ix10234 : nand03 port map ( Y=>nx10233, A0=>nx14440, A1=>nx2484, A2=>
      nx14434);
   ix2485 : xnor2 port map ( Y=>nx2484, A0=>nx2328, A1=>nx10246);
   ix2329 : oai22 port map ( Y=>nx2328, A0=>nx10217, A1=>nx10227, B0=>
      nx10231, B1=>nx10237);
   ix10245 : inv01 port map ( Y=>nx10244, A=>weight_7(10));
   ix10247 : xnor2 port map ( Y=>nx10246, A0=>
      booth_integrtaion_7_booth_output_27, A1=>nx2348);
   booth_integrtaion_7_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_27, QB=>OPEN, D=>nx4331, CLK=>clk, R
      =>rst);
   ix10252 : xnor2 port map ( Y=>nx10251, A0=>nx10253, A1=>nx10263);
   ix10254 : aoi22 port map ( Y=>nx10253, A0=>
      booth_integrtaion_7_booth_output_27, A1=>nx2348, B0=>nx2328, B1=>
      nx2881);
   ix2349 : oai32 port map ( Y=>nx2348, A0=>nx10256, A1=>nx14446, A2=>nx2338, 
      B0=>nx10260, B1=>nx14450);
   ix10257 : nor02ii port map ( Y=>nx10256, A0=>nx2314, A1=>weight_7(11));
   ix2315 : nor02ii port map ( Y=>nx2314, A0=>weight_7(10), A1=>nx2290);
   ix2339 : nor02ii port map ( Y=>nx2338, A0=>weight_7(11), A1=>nx2314);
   ix10261 : inv01 port map ( Y=>nx10260, A=>weight_7(11));
   ix4322 : oai21 port map ( Y=>nx4321, A0=>nx10267, A1=>nx14434, B0=>
      nx10269);
   booth_integrtaion_7_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10267, D=>nx4321, CLK=>clk, R=>rst);
   ix10270 : nand03 port map ( Y=>nx10269, A0=>nx14698, A1=>nx2460, A2=>
      nx14434);
   ix2461 : xnor2 port map ( Y=>nx2460, A0=>nx2376, A1=>nx10282);
   ix2377 : oai22 port map ( Y=>nx2376, A0=>nx10253, A1=>nx10263, B0=>
      nx10267, B1=>nx10273);
   ix10281 : inv01 port map ( Y=>nx10280, A=>weight_7(12));
   ix10283 : xnor2 port map ( Y=>nx10282, A0=>
      booth_integrtaion_7_booth_output_29, A1=>nx2396);
   booth_integrtaion_7_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_29, QB=>OPEN, D=>nx4311, CLK=>clk, R
      =>rst);
   ix10288 : xnor2 port map ( Y=>nx10287, A0=>nx10289, A1=>nx10299);
   ix10290 : aoi22 port map ( Y=>nx10289, A0=>
      booth_integrtaion_7_booth_output_29, A1=>nx2396, B0=>nx2376, B1=>
      nx2885);
   ix2397 : oai32 port map ( Y=>nx2396, A0=>nx10292, A1=>nx14446, A2=>nx2386, 
      B0=>nx10296, B1=>nx14450);
   ix10293 : nor02ii port map ( Y=>nx10292, A0=>nx2362, A1=>weight_7(13));
   ix2363 : nor02ii port map ( Y=>nx2362, A0=>weight_7(12), A1=>nx2338);
   ix2387 : nor02ii port map ( Y=>nx2386, A0=>weight_7(13), A1=>nx2362);
   ix10297 : inv01 port map ( Y=>nx10296, A=>weight_7(13));
   ix10305 : xnor2 port map ( Y=>nx10304, A0=>nx2424, A1=>nx2434);
   ix2425 : oai22 port map ( Y=>nx2424, A0=>nx10289, A1=>nx10299, B0=>
      nx10307, B1=>nx10309);
   booth_integrtaion_7_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_31, QB=>nx10307, D=>nx4301, CLK=>clk, 
      R=>rst);
   ix10317 : inv01 port map ( Y=>nx10316, A=>weight_7(14));
   ix10320 : aoi22 port map ( Y=>nx10319, A0=>weight_7(15), A1=>nx2074, B0=>
      nx2078, B1=>nx2426);
   ix2427 : xnor2 port map ( Y=>nx2426, A0=>weight_7(15), A1=>nx2410);
   ix2411 : nor02ii port map ( Y=>nx2410, A0=>weight_7(14), A1=>nx2386);
   ix2421 : oai32 port map ( Y=>nx2420, A0=>nx10324, A1=>nx14446, A2=>nx2410, 
      B0=>nx10316, B1=>nx14450);
   ix10325 : nor02ii port map ( Y=>nx10324, A0=>nx2386, A1=>weight_7(14));
   ix2373 : oai32 port map ( Y=>nx2372, A0=>nx10328, A1=>nx14448, A2=>nx2362, 
      B0=>nx10280, B1=>nx14452);
   ix10329 : nor02ii port map ( Y=>nx10328, A0=>nx2338, A1=>weight_7(12));
   ix2325 : oai32 port map ( Y=>nx2324, A0=>nx10332, A1=>nx14448, A2=>nx2314, 
      B0=>nx10244, B1=>nx14452);
   ix10333 : nor02ii port map ( Y=>nx10332, A0=>nx2290, A1=>weight_7(10));
   ix2277 : oai32 port map ( Y=>nx2276, A0=>nx10336, A1=>nx14448, A2=>nx2266, 
      B0=>nx10208, B1=>nx14452);
   ix10337 : nor02ii port map ( Y=>nx10336, A0=>nx2242, A1=>weight_7(8));
   ix2229 : oai32 port map ( Y=>nx2228, A0=>nx10340, A1=>nx14448, A2=>nx2218, 
      B0=>nx10172, B1=>nx14452);
   ix10341 : nor02ii port map ( Y=>nx10340, A0=>nx2194, A1=>weight_7(6));
   ix2181 : oai32 port map ( Y=>nx2180, A0=>nx10344, A1=>nx14448, A2=>nx2170, 
      B0=>nx10136, B1=>nx14452);
   ix10345 : nor02ii port map ( Y=>nx10344, A0=>nx2146, A1=>weight_7(4));
   ix10348 : aoi32 port map ( Y=>nx10347, A0=>nx2092, A1=>nx2078, A2=>
      nx10080, B0=>weight_7(1), B1=>nx2074);
   booth_integrtaion_7_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_7_booth_output_16, QB=>nx10061, D=>nx4441, CLK=>clk, 
      R=>rst);
   booth_integrtaion_7_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_7_15, QB=>nx10351, D=>nx4451, CLK=>clk, R=>
      rst);
   ix2957 : xor2 port map ( Y=>label_7(1), A0=>nx10368, A1=>nx10370);
   ix10369 : nand02 port map ( Y=>nx10368, A0=>adderInput_7(0), A1=>
      booth_integration_output_7_0);
   ix10371 : xnor2 port map ( Y=>nx10370, A0=>booth_integration_output_7_1, 
      A1=>adderInput_7(1));
   ix2955 : xor2 port map ( Y=>label_7(2), A0=>nx10373, A1=>nx10376);
   ix10374 : aoi32 port map ( Y=>nx10373, A0=>adderInput_7(0), A1=>
      booth_integration_output_7_0, A2=>nx2814, B0=>adderInput_7(1), B1=>
      booth_integration_output_7_1);
   ix2953 : xnor2 port map ( Y=>label_7(3), A0=>nx2828, A1=>nx10382);
   ix2829 : oai22 port map ( Y=>nx2828, A0=>nx10373, A1=>nx10376, B0=>
      nx10380, B1=>nx10365);
   ix10381 : inv01 port map ( Y=>nx10380, A=>adderInput_7(2));
   ix10383 : xnor2 port map ( Y=>nx10382, A0=>booth_integration_output_7_3, 
      A1=>adderInput_7(3));
   ix2951 : xor2 port map ( Y=>label_7(4), A0=>nx10385, A1=>nx10388);
   ix10386 : aoi22 port map ( Y=>nx10385, A0=>adderInput_7(3), A1=>
      booth_integration_output_7_3, B0=>nx2828, B1=>nx2830);
   ix2949 : xnor2 port map ( Y=>label_7(5), A0=>nx2844, A1=>nx10394);
   ix2845 : oai22 port map ( Y=>nx2844, A0=>nx10385, A1=>nx10388, B0=>
      nx10392, B1=>nx10363);
   ix10393 : inv01 port map ( Y=>nx10392, A=>adderInput_7(4));
   ix10395 : xnor2 port map ( Y=>nx10394, A0=>booth_integration_output_7_5, 
      A1=>adderInput_7(5));
   ix2947 : xor2 port map ( Y=>label_7(6), A0=>nx10397, A1=>nx10400);
   ix10398 : aoi22 port map ( Y=>nx10397, A0=>adderInput_7(5), A1=>
      booth_integration_output_7_5, B0=>nx2844, B1=>nx2846);
   ix2945 : xnor2 port map ( Y=>label_7(7), A0=>nx2860, A1=>nx10406);
   ix2861 : oai22 port map ( Y=>nx2860, A0=>nx10397, A1=>nx10400, B0=>
      nx10404, B1=>nx10361);
   ix10405 : inv01 port map ( Y=>nx10404, A=>adderInput_7(6));
   ix10407 : xnor2 port map ( Y=>nx10406, A0=>booth_integration_output_7_7, 
      A1=>adderInput_7(7));
   ix2943 : xor2 port map ( Y=>label_7(8), A0=>nx10409, A1=>nx10412);
   ix10410 : aoi22 port map ( Y=>nx10409, A0=>adderInput_7(7), A1=>
      booth_integration_output_7_7, B0=>nx2860, B1=>nx2862);
   ix2941 : xnor2 port map ( Y=>label_7(9), A0=>nx2876, A1=>nx10418);
   ix2877 : oai22 port map ( Y=>nx2876, A0=>nx10409, A1=>nx10412, B0=>
      nx10416, B1=>nx10359);
   ix10417 : inv01 port map ( Y=>nx10416, A=>adderInput_7(8));
   ix10419 : xnor2 port map ( Y=>nx10418, A0=>booth_integration_output_7_9, 
      A1=>adderInput_7(9));
   ix2939 : xor2 port map ( Y=>label_7(10), A0=>nx10421, A1=>nx10424);
   ix10422 : aoi22 port map ( Y=>nx10421, A0=>adderInput_7(9), A1=>
      booth_integration_output_7_9, B0=>nx2876, B1=>nx2878);
   ix2937 : xnor2 port map ( Y=>label_7(11), A0=>nx2892, A1=>nx10430);
   ix2893 : oai22 port map ( Y=>nx2892, A0=>nx10421, A1=>nx10424, B0=>
      nx10428, B1=>nx10357);
   ix10429 : inv01 port map ( Y=>nx10428, A=>adderInput_7(10));
   ix10431 : xnor2 port map ( Y=>nx10430, A0=>booth_integration_output_7_11, 
      A1=>adderInput_7(11));
   ix2935 : xor2 port map ( Y=>label_7(12), A0=>nx10433, A1=>nx10436);
   ix10434 : aoi22 port map ( Y=>nx10433, A0=>adderInput_7(11), A1=>
      booth_integration_output_7_11, B0=>nx2892, B1=>nx2894);
   ix2933 : xnor2 port map ( Y=>label_7(13), A0=>nx2908, A1=>nx10442);
   ix2909 : oai22 port map ( Y=>nx2908, A0=>nx10433, A1=>nx10436, B0=>
      nx10440, B1=>nx10355);
   ix10441 : inv01 port map ( Y=>nx10440, A=>adderInput_7(12));
   ix10443 : xnor2 port map ( Y=>nx10442, A0=>booth_integration_output_7_13, 
      A1=>adderInput_7(13));
   ix2931 : xor2 port map ( Y=>label_7(14), A0=>nx10445, A1=>nx10448);
   ix10446 : aoi22 port map ( Y=>nx10445, A0=>adderInput_7(13), A1=>
      booth_integration_output_7_13, B0=>nx2908, B1=>nx2910);
   ix2929 : xnor2 port map ( Y=>label_7(15), A0=>nx2924, A1=>nx10454);
   ix2925 : oai22 port map ( Y=>nx2924, A0=>nx10445, A1=>nx10448, B0=>
      nx10452, B1=>nx10353);
   ix10453 : inv01 port map ( Y=>nx10452, A=>adderInput_7(14));
   booth_integrtaion_6_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_1, QB=>OPEN, D=>nx5121, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_2, QB=>nx10888, D=>nx5111, CLK=>clk, R=>rst
   );
   booth_integrtaion_6_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_3, QB=>OPEN, D=>nx5101, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_4, QB=>nx10886, D=>nx5091, CLK=>clk, R=>rst
   );
   booth_integrtaion_6_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_5, QB=>OPEN, D=>nx5081, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_6, QB=>nx10884, D=>nx5071, CLK=>clk, R=>rst
   );
   booth_integrtaion_6_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_7, QB=>OPEN, D=>nx5061, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_8, QB=>nx10882, D=>nx5051, CLK=>clk, R=>rst
   );
   booth_integrtaion_6_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_9, QB=>OPEN, D=>nx5041, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_10, QB=>nx10880, D=>nx5031, CLK=>clk, R=>
      rst);
   booth_integrtaion_6_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_11, QB=>OPEN, D=>nx5021, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_12, QB=>nx10878, D=>nx5011, CLK=>clk, R=>
      rst);
   booth_integrtaion_6_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_13, QB=>OPEN, D=>nx5001, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_14, QB=>nx10876, D=>nx4991, CLK=>clk, R=>
      rst);
   ix10506 : aoi22 port map ( Y=>nx10505, A0=>neuron(15), A1=>nx14240, B0=>
      nx3600, B1=>nx3606);
   booth_integrtaion_6_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_reg_output_0, QB=>OPEN, D=>nx4631, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_0, QB=>OPEN, D=>nx4617, CLK=>clk, 
      S=>nx14154);
   booth_integrtaion_6_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_reg_output_9, QB=>OPEN, D=>nx4811, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_9, QB=>OPEN, D=>nx4801, CLK=>clk, 
      R=>nx14152);
   booth_integrtaion_6_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_8, QB=>OPEN, D=>nx4791, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_8, QB=>OPEN, D=>nx4781, CLK=>clk, 
      R=>nx14152);
   booth_integrtaion_6_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_7, QB=>OPEN, D=>nx4771, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_7, QB=>OPEN, D=>nx4761, CLK=>clk, 
      R=>nx14152);
   booth_integrtaion_6_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_6, QB=>OPEN, D=>nx4751, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_6, QB=>OPEN, D=>nx4741, CLK=>clk, 
      R=>nx14152);
   booth_integrtaion_6_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_5, QB=>OPEN, D=>nx4731, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_5, QB=>OPEN, D=>nx4721, CLK=>clk, 
      R=>nx14152);
   booth_integrtaion_6_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_4, QB=>OPEN, D=>nx4711, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_4, QB=>OPEN, D=>nx4701, CLK=>clk, 
      R=>nx14152);
   booth_integrtaion_6_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_3, QB=>OPEN, D=>nx4691, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_3, QB=>OPEN, D=>nx4681, CLK=>clk, 
      R=>nx14152);
   booth_integrtaion_6_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_2, QB=>OPEN, D=>nx4671, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_2, QB=>OPEN, D=>nx4661, CLK=>clk, 
      R=>nx14150);
   booth_integrtaion_6_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_output_1, QB=>OPEN, D=>nx4651, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_6_shift_Reg_count_1, QB=>OPEN, D=>nx4641, CLK=>clk, 
      R=>nx14150);
   ix4612 : nand02 port map ( Y=>nx4611, A0=>nx14624, A1=>nx14226);
   booth_integrtaion_6_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx10552, D=>nx4611, CLK=>clk, S=>nx14150);
   ix3601 : nand02 port map ( Y=>nx3600, A0=>nx10573, A1=>nx10584);
   ix10574 : oai21 port map ( Y=>nx10573, A0=>nx3064, A1=>nx3060, B0=>
      weight_6(0));
   ix4822 : oai21 port map ( Y=>nx4821, A0=>nx10578, A1=>nx14454, B0=>
      nx10580);
   booth_integrtaion_6_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10578, D=>nx4821, CLK=>clk, R=>rst);
   booth_integrtaion_6_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_0, QB=>nx10457, D=>nx5131, CLK=>clk, R=>rst
   );
   ix10589 : xnor2 port map ( Y=>nx10588, A0=>nx3070, A1=>nx2891);
   ix4962 : oai21 port map ( Y=>nx4961, A0=>nx10594, A1=>nx14454, B0=>
      nx10596);
   booth_integrtaion_6_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_17, QB=>nx10594, D=>nx4961, CLK=>clk, 
      R=>rst);
   ix10597 : nand03 port map ( Y=>nx10596, A0=>nx14462, A1=>nx3578, A2=>
      nx14706);
   ix3579 : xnor2 port map ( Y=>nx3578, A0=>nx10599, A1=>nx2893);
   ix10600 : aoi22 port map ( Y=>nx10599, A0=>
      booth_integrtaion_6_booth_output_17, A1=>nx3094, B0=>nx3070, B1=>
      nx2891);
   ix3079 : nand02 port map ( Y=>nx3078, A0=>weight_6(1), A1=>weight_6(0));
   ix10604 : or02 port map ( Y=>nx10603, A0=>weight_6(0), A1=>weight_6(1));
   ix4952 : oai21 port map ( Y=>nx4951, A0=>nx10608, A1=>nx14454, B0=>
      nx10610);
   booth_integrtaion_6_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10608, D=>nx4951, CLK=>clk, R=>rst);
   ix10611 : nand03 port map ( Y=>nx10610, A0=>nx14462, A1=>nx3566, A2=>
      nx14706);
   ix3567 : xnor2 port map ( Y=>nx3566, A0=>nx3122, A1=>nx10621);
   ix3123 : oai22 port map ( Y=>nx3122, A0=>nx10599, A1=>nx10614, B0=>
      nx10608, B1=>nx14466);
   ix10617 : aoi32 port map ( Y=>nx10616, A0=>nx3104, A1=>nx3064, A2=>
      nx10619, B0=>weight_6(2), B1=>nx3060);
   ix3105 : oai21 port map ( Y=>nx3104, A0=>weight_6(0), A1=>weight_6(1), B0
      =>weight_6(2));
   ix10622 : xnor2 port map ( Y=>nx10621, A0=>
      booth_integrtaion_6_booth_output_19, A1=>nx3142);
   booth_integrtaion_6_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_19, QB=>OPEN, D=>nx4941, CLK=>clk, R
      =>rst);
   ix10627 : xnor2 port map ( Y=>nx10626, A0=>nx10628, A1=>nx10642);
   ix10629 : aoi22 port map ( Y=>nx10628, A0=>
      booth_integrtaion_6_booth_output_19, A1=>nx3142, B0=>nx3122, B1=>
      nx2895);
   ix3143 : oai32 port map ( Y=>nx3142, A0=>nx10631, A1=>nx14468, A2=>nx3132, 
      B0=>nx10637, B1=>nx14472);
   ix10632 : nor02ii port map ( Y=>nx10631, A0=>nx3108, A1=>weight_6(3));
   ix3109 : nor03_2x port map ( Y=>nx3108, A0=>weight_6(2), A1=>weight_6(0), 
      A2=>weight_6(1));
   ix3133 : nor04 port map ( Y=>nx3132, A0=>weight_6(3), A1=>weight_6(2), A2
      =>weight_6(0), A3=>weight_6(1));
   ix10638 : inv01 port map ( Y=>nx10637, A=>weight_6(3));
   ix4932 : oai21 port map ( Y=>nx4931, A0=>nx10646, A1=>nx14454, B0=>
      nx10648);
   booth_integrtaion_6_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10646, D=>nx4931, CLK=>clk, R=>rst);
   ix10649 : nand03 port map ( Y=>nx10648, A0=>nx14462, A1=>nx3542, A2=>
      nx14706);
   ix3543 : xnor2 port map ( Y=>nx3542, A0=>nx3170, A1=>nx10661);
   ix3171 : oai22 port map ( Y=>nx3170, A0=>nx10628, A1=>nx10642, B0=>
      nx10646, B1=>nx10652);
   ix10660 : inv01 port map ( Y=>nx10659, A=>weight_6(4));
   ix10662 : xnor2 port map ( Y=>nx10661, A0=>
      booth_integrtaion_6_booth_output_21, A1=>nx3190);
   booth_integrtaion_6_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_21, QB=>OPEN, D=>nx4921, CLK=>clk, R
      =>rst);
   ix10667 : xnor2 port map ( Y=>nx10666, A0=>nx10668, A1=>nx10678);
   ix10669 : aoi22 port map ( Y=>nx10668, A0=>
      booth_integrtaion_6_booth_output_21, A1=>nx3190, B0=>nx3170, B1=>
      nx2899);
   ix3191 : oai32 port map ( Y=>nx3190, A0=>nx10671, A1=>nx14468, A2=>nx3180, 
      B0=>nx10675, B1=>nx14472);
   ix10672 : nor02ii port map ( Y=>nx10671, A0=>nx3156, A1=>weight_6(5));
   ix3157 : nor02ii port map ( Y=>nx3156, A0=>weight_6(4), A1=>nx3132);
   ix3181 : nor02ii port map ( Y=>nx3180, A0=>weight_6(5), A1=>nx3156);
   ix10676 : inv01 port map ( Y=>nx10675, A=>weight_6(5));
   ix4912 : oai21 port map ( Y=>nx4911, A0=>nx10682, A1=>nx14454, B0=>
      nx10684);
   booth_integrtaion_6_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10682, D=>nx4911, CLK=>clk, R=>rst);
   ix10685 : nand03 port map ( Y=>nx10684, A0=>nx14462, A1=>nx3518, A2=>
      nx14456);
   ix3519 : xnor2 port map ( Y=>nx3518, A0=>nx3218, A1=>nx10697);
   ix3219 : oai22 port map ( Y=>nx3218, A0=>nx10668, A1=>nx10678, B0=>
      nx10682, B1=>nx10688);
   ix10696 : inv01 port map ( Y=>nx10695, A=>weight_6(6));
   ix10698 : xnor2 port map ( Y=>nx10697, A0=>
      booth_integrtaion_6_booth_output_23, A1=>nx3238);
   booth_integrtaion_6_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_23, QB=>OPEN, D=>nx4901, CLK=>clk, R
      =>rst);
   ix10703 : xnor2 port map ( Y=>nx10702, A0=>nx10704, A1=>nx10714);
   ix10705 : aoi22 port map ( Y=>nx10704, A0=>
      booth_integrtaion_6_booth_output_23, A1=>nx3238, B0=>nx3218, B1=>
      nx2903);
   ix3239 : oai32 port map ( Y=>nx3238, A0=>nx10707, A1=>nx14468, A2=>nx3228, 
      B0=>nx10711, B1=>nx14472);
   ix10708 : nor02ii port map ( Y=>nx10707, A0=>nx3204, A1=>weight_6(7));
   ix3205 : nor02ii port map ( Y=>nx3204, A0=>weight_6(6), A1=>nx3180);
   ix3229 : nor02ii port map ( Y=>nx3228, A0=>weight_6(7), A1=>nx3204);
   ix10712 : inv01 port map ( Y=>nx10711, A=>weight_6(7));
   ix4892 : oai21 port map ( Y=>nx4891, A0=>nx10718, A1=>nx14456, B0=>
      nx10720);
   booth_integrtaion_6_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10718, D=>nx4891, CLK=>clk, R=>rst);
   ix10721 : nand03 port map ( Y=>nx10720, A0=>nx14462, A1=>nx3494, A2=>
      nx14456);
   ix3495 : xnor2 port map ( Y=>nx3494, A0=>nx3266, A1=>nx10733);
   ix3267 : oai22 port map ( Y=>nx3266, A0=>nx10704, A1=>nx10714, B0=>
      nx10718, B1=>nx10724);
   ix10732 : inv01 port map ( Y=>nx10731, A=>weight_6(8));
   ix10734 : xnor2 port map ( Y=>nx10733, A0=>
      booth_integrtaion_6_booth_output_25, A1=>nx3286);
   booth_integrtaion_6_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_25, QB=>OPEN, D=>nx4881, CLK=>clk, R
      =>rst);
   ix10739 : xnor2 port map ( Y=>nx10738, A0=>nx10740, A1=>nx10750);
   ix10741 : aoi22 port map ( Y=>nx10740, A0=>
      booth_integrtaion_6_booth_output_25, A1=>nx3286, B0=>nx3266, B1=>
      nx2907);
   ix3287 : oai32 port map ( Y=>nx3286, A0=>nx10743, A1=>nx14468, A2=>nx3276, 
      B0=>nx10747, B1=>nx14472);
   ix10744 : nor02ii port map ( Y=>nx10743, A0=>nx3252, A1=>weight_6(9));
   ix3253 : nor02ii port map ( Y=>nx3252, A0=>weight_6(8), A1=>nx3228);
   ix3277 : nor02ii port map ( Y=>nx3276, A0=>weight_6(9), A1=>nx3252);
   ix10748 : inv01 port map ( Y=>nx10747, A=>weight_6(9));
   ix4872 : oai21 port map ( Y=>nx4871, A0=>nx10754, A1=>nx14456, B0=>
      nx10756);
   booth_integrtaion_6_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10754, D=>nx4871, CLK=>clk, R=>rst);
   ix10757 : nand03 port map ( Y=>nx10756, A0=>nx14462, A1=>nx3470, A2=>
      nx14456);
   ix3471 : xnor2 port map ( Y=>nx3470, A0=>nx3314, A1=>nx10769);
   ix3315 : oai22 port map ( Y=>nx3314, A0=>nx10740, A1=>nx10750, B0=>
      nx10754, B1=>nx10760);
   ix10768 : inv01 port map ( Y=>nx10767, A=>weight_6(10));
   ix10770 : xnor2 port map ( Y=>nx10769, A0=>
      booth_integrtaion_6_booth_output_27, A1=>nx3334);
   booth_integrtaion_6_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_27, QB=>OPEN, D=>nx4861, CLK=>clk, R
      =>rst);
   ix10775 : xnor2 port map ( Y=>nx10774, A0=>nx10776, A1=>nx10786);
   ix10777 : aoi22 port map ( Y=>nx10776, A0=>
      booth_integrtaion_6_booth_output_27, A1=>nx3334, B0=>nx3314, B1=>
      nx2911);
   ix3335 : oai32 port map ( Y=>nx3334, A0=>nx10779, A1=>nx14468, A2=>nx3324, 
      B0=>nx10783, B1=>nx14472);
   ix10780 : nor02ii port map ( Y=>nx10779, A0=>nx3300, A1=>weight_6(11));
   ix3301 : nor02ii port map ( Y=>nx3300, A0=>weight_6(10), A1=>nx3276);
   ix3325 : nor02ii port map ( Y=>nx3324, A0=>weight_6(11), A1=>nx3300);
   ix10784 : inv01 port map ( Y=>nx10783, A=>weight_6(11));
   ix4852 : oai21 port map ( Y=>nx4851, A0=>nx10790, A1=>nx14456, B0=>
      nx10792);
   booth_integrtaion_6_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx10790, D=>nx4851, CLK=>clk, R=>rst);
   ix10793 : nand03 port map ( Y=>nx10792, A0=>nx14714, A1=>nx3446, A2=>
      nx14456);
   ix3447 : xnor2 port map ( Y=>nx3446, A0=>nx3362, A1=>nx10805);
   ix3363 : oai22 port map ( Y=>nx3362, A0=>nx10776, A1=>nx10786, B0=>
      nx10790, B1=>nx10796);
   ix10804 : inv01 port map ( Y=>nx10803, A=>weight_6(12));
   ix10806 : xnor2 port map ( Y=>nx10805, A0=>
      booth_integrtaion_6_booth_output_29, A1=>nx3382);
   booth_integrtaion_6_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_29, QB=>OPEN, D=>nx4841, CLK=>clk, R
      =>rst);
   ix10811 : xnor2 port map ( Y=>nx10810, A0=>nx10812, A1=>nx10822);
   ix10813 : aoi22 port map ( Y=>nx10812, A0=>
      booth_integrtaion_6_booth_output_29, A1=>nx3382, B0=>nx3362, B1=>
      nx2915);
   ix3383 : oai32 port map ( Y=>nx3382, A0=>nx10815, A1=>nx14468, A2=>nx3372, 
      B0=>nx10819, B1=>nx14472);
   ix10816 : nor02ii port map ( Y=>nx10815, A0=>nx3348, A1=>weight_6(13));
   ix3349 : nor02ii port map ( Y=>nx3348, A0=>weight_6(12), A1=>nx3324);
   ix3373 : nor02ii port map ( Y=>nx3372, A0=>weight_6(13), A1=>nx3348);
   ix10820 : inv01 port map ( Y=>nx10819, A=>weight_6(13));
   ix10828 : xnor2 port map ( Y=>nx10827, A0=>nx3410, A1=>nx3420);
   ix3411 : oai22 port map ( Y=>nx3410, A0=>nx10812, A1=>nx10822, B0=>
      nx10830, B1=>nx10832);
   booth_integrtaion_6_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_31, QB=>nx10830, D=>nx4831, CLK=>clk, 
      R=>rst);
   ix10840 : inv01 port map ( Y=>nx10839, A=>weight_6(14));
   ix10843 : aoi22 port map ( Y=>nx10842, A0=>weight_6(15), A1=>nx3060, B0=>
      nx3064, B1=>nx3412);
   ix3413 : xnor2 port map ( Y=>nx3412, A0=>weight_6(15), A1=>nx3396);
   ix3397 : nor02ii port map ( Y=>nx3396, A0=>weight_6(14), A1=>nx3372);
   ix3407 : oai32 port map ( Y=>nx3406, A0=>nx10847, A1=>nx14468, A2=>nx3396, 
      B0=>nx10839, B1=>nx14472);
   ix10848 : nor02ii port map ( Y=>nx10847, A0=>nx3372, A1=>weight_6(14));
   ix3359 : oai32 port map ( Y=>nx3358, A0=>nx10851, A1=>nx14470, A2=>nx3348, 
      B0=>nx10803, B1=>nx14474);
   ix10852 : nor02ii port map ( Y=>nx10851, A0=>nx3324, A1=>weight_6(12));
   ix3311 : oai32 port map ( Y=>nx3310, A0=>nx10855, A1=>nx14470, A2=>nx3300, 
      B0=>nx10767, B1=>nx14474);
   ix10856 : nor02ii port map ( Y=>nx10855, A0=>nx3276, A1=>weight_6(10));
   ix3263 : oai32 port map ( Y=>nx3262, A0=>nx10859, A1=>nx14470, A2=>nx3252, 
      B0=>nx10731, B1=>nx14474);
   ix10860 : nor02ii port map ( Y=>nx10859, A0=>nx3228, A1=>weight_6(8));
   ix3215 : oai32 port map ( Y=>nx3214, A0=>nx10863, A1=>nx14470, A2=>nx3204, 
      B0=>nx10695, B1=>nx14474);
   ix10864 : nor02ii port map ( Y=>nx10863, A0=>nx3180, A1=>weight_6(6));
   ix3167 : oai32 port map ( Y=>nx3166, A0=>nx10867, A1=>nx14470, A2=>nx3156, 
      B0=>nx10659, B1=>nx14474);
   ix10868 : nor02ii port map ( Y=>nx10867, A0=>nx3132, A1=>weight_6(4));
   ix10871 : aoi32 port map ( Y=>nx10870, A0=>nx3078, A1=>nx3064, A2=>
      nx10603, B0=>weight_6(1), B1=>nx3060);
   booth_integrtaion_6_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_6_booth_output_16, QB=>nx10584, D=>nx4971, CLK=>clk, 
      R=>rst);
   booth_integrtaion_6_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_6_15, QB=>nx10874, D=>nx4981, CLK=>clk, R=>
      rst);
   ix3943 : xor2 port map ( Y=>label_6(1), A0=>nx10891, A1=>nx10893);
   ix10892 : nand02 port map ( Y=>nx10891, A0=>adderInput_6(0), A1=>
      booth_integration_output_6_0);
   ix10894 : xnor2 port map ( Y=>nx10893, A0=>booth_integration_output_6_1, 
      A1=>adderInput_6(1));
   ix3941 : xor2 port map ( Y=>label_6(2), A0=>nx10896, A1=>nx10899);
   ix10897 : aoi32 port map ( Y=>nx10896, A0=>adderInput_6(0), A1=>
      booth_integration_output_6_0, A2=>nx3800, B0=>adderInput_6(1), B1=>
      booth_integration_output_6_1);
   ix3939 : xnor2 port map ( Y=>label_6(3), A0=>nx3814, A1=>nx10905);
   ix3815 : oai22 port map ( Y=>nx3814, A0=>nx10896, A1=>nx10899, B0=>
      nx10903, B1=>nx10888);
   ix10904 : inv01 port map ( Y=>nx10903, A=>adderInput_6(2));
   ix10906 : xnor2 port map ( Y=>nx10905, A0=>booth_integration_output_6_3, 
      A1=>adderInput_6(3));
   ix3937 : xor2 port map ( Y=>label_6(4), A0=>nx10908, A1=>nx10911);
   ix10909 : aoi22 port map ( Y=>nx10908, A0=>adderInput_6(3), A1=>
      booth_integration_output_6_3, B0=>nx3814, B1=>nx3816);
   ix3935 : xnor2 port map ( Y=>label_6(5), A0=>nx3830, A1=>nx10917);
   ix3831 : oai22 port map ( Y=>nx3830, A0=>nx10908, A1=>nx10911, B0=>
      nx10915, B1=>nx10886);
   ix10916 : inv01 port map ( Y=>nx10915, A=>adderInput_6(4));
   ix10918 : xnor2 port map ( Y=>nx10917, A0=>booth_integration_output_6_5, 
      A1=>adderInput_6(5));
   ix3933 : xor2 port map ( Y=>label_6(6), A0=>nx10920, A1=>nx10923);
   ix10921 : aoi22 port map ( Y=>nx10920, A0=>adderInput_6(5), A1=>
      booth_integration_output_6_5, B0=>nx3830, B1=>nx3832);
   ix3931 : xnor2 port map ( Y=>label_6(7), A0=>nx3846, A1=>nx10929);
   ix3847 : oai22 port map ( Y=>nx3846, A0=>nx10920, A1=>nx10923, B0=>
      nx10927, B1=>nx10884);
   ix10928 : inv01 port map ( Y=>nx10927, A=>adderInput_6(6));
   ix10930 : xnor2 port map ( Y=>nx10929, A0=>booth_integration_output_6_7, 
      A1=>adderInput_6(7));
   ix3929 : xor2 port map ( Y=>label_6(8), A0=>nx10932, A1=>nx10935);
   ix10933 : aoi22 port map ( Y=>nx10932, A0=>adderInput_6(7), A1=>
      booth_integration_output_6_7, B0=>nx3846, B1=>nx3848);
   ix3927 : xnor2 port map ( Y=>label_6(9), A0=>nx3862, A1=>nx10941);
   ix3863 : oai22 port map ( Y=>nx3862, A0=>nx10932, A1=>nx10935, B0=>
      nx10939, B1=>nx10882);
   ix10940 : inv01 port map ( Y=>nx10939, A=>adderInput_6(8));
   ix10942 : xnor2 port map ( Y=>nx10941, A0=>booth_integration_output_6_9, 
      A1=>adderInput_6(9));
   ix3925 : xor2 port map ( Y=>label_6(10), A0=>nx10944, A1=>nx10947);
   ix10945 : aoi22 port map ( Y=>nx10944, A0=>adderInput_6(9), A1=>
      booth_integration_output_6_9, B0=>nx3862, B1=>nx3864);
   ix3923 : xnor2 port map ( Y=>label_6(11), A0=>nx3878, A1=>nx10953);
   ix3879 : oai22 port map ( Y=>nx3878, A0=>nx10944, A1=>nx10947, B0=>
      nx10951, B1=>nx10880);
   ix10952 : inv01 port map ( Y=>nx10951, A=>adderInput_6(10));
   ix10954 : xnor2 port map ( Y=>nx10953, A0=>booth_integration_output_6_11, 
      A1=>adderInput_6(11));
   ix3921 : xor2 port map ( Y=>label_6(12), A0=>nx10956, A1=>nx10959);
   ix10957 : aoi22 port map ( Y=>nx10956, A0=>adderInput_6(11), A1=>
      booth_integration_output_6_11, B0=>nx3878, B1=>nx3880);
   ix3919 : xnor2 port map ( Y=>label_6(13), A0=>nx3894, A1=>nx10965);
   ix3895 : oai22 port map ( Y=>nx3894, A0=>nx10956, A1=>nx10959, B0=>
      nx10963, B1=>nx10878);
   ix10964 : inv01 port map ( Y=>nx10963, A=>adderInput_6(12));
   ix10966 : xnor2 port map ( Y=>nx10965, A0=>booth_integration_output_6_13, 
      A1=>adderInput_6(13));
   ix3917 : xor2 port map ( Y=>label_6(14), A0=>nx10968, A1=>nx10971);
   ix10969 : aoi22 port map ( Y=>nx10968, A0=>adderInput_6(13), A1=>
      booth_integration_output_6_13, B0=>nx3894, B1=>nx3896);
   ix3915 : xnor2 port map ( Y=>label_6(15), A0=>nx3910, A1=>nx10977);
   ix3911 : oai22 port map ( Y=>nx3910, A0=>nx10968, A1=>nx10971, B0=>
      nx10975, B1=>nx10876);
   ix10976 : inv01 port map ( Y=>nx10975, A=>adderInput_6(14));
   booth_integrtaion_5_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_1, QB=>OPEN, D=>nx5651, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_2, QB=>nx11411, D=>nx5641, CLK=>clk, R=>rst
   );
   booth_integrtaion_5_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_3, QB=>OPEN, D=>nx5631, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_4, QB=>nx11409, D=>nx5621, CLK=>clk, R=>rst
   );
   booth_integrtaion_5_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_5, QB=>OPEN, D=>nx5611, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_6, QB=>nx11407, D=>nx5601, CLK=>clk, R=>rst
   );
   booth_integrtaion_5_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_7, QB=>OPEN, D=>nx5591, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_8, QB=>nx11405, D=>nx5581, CLK=>clk, R=>rst
   );
   booth_integrtaion_5_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_9, QB=>OPEN, D=>nx5571, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_10, QB=>nx11403, D=>nx5561, CLK=>clk, R=>
      rst);
   booth_integrtaion_5_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_11, QB=>OPEN, D=>nx5551, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_12, QB=>nx11401, D=>nx5541, CLK=>clk, R=>
      rst);
   booth_integrtaion_5_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_13, QB=>OPEN, D=>nx5531, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_14, QB=>nx11399, D=>nx5521, CLK=>clk, R=>
      rst);
   ix11029 : aoi22 port map ( Y=>nx11028, A0=>neuron(15), A1=>nx14262, B0=>
      nx4586, B1=>nx4592);
   booth_integrtaion_5_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_reg_output_0, QB=>OPEN, D=>nx5161, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_0, QB=>OPEN, D=>nx5147, CLK=>clk, 
      S=>nx14156);
   booth_integrtaion_5_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_reg_output_9, QB=>OPEN, D=>nx5341, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_9, QB=>OPEN, D=>nx5331, CLK=>clk, 
      R=>nx14156);
   booth_integrtaion_5_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_8, QB=>OPEN, D=>nx5321, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_8, QB=>OPEN, D=>nx5311, CLK=>clk, 
      R=>nx14156);
   booth_integrtaion_5_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_7, QB=>OPEN, D=>nx5301, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_7, QB=>OPEN, D=>nx5291, CLK=>clk, 
      R=>nx14156);
   booth_integrtaion_5_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_6, QB=>OPEN, D=>nx5281, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_6, QB=>OPEN, D=>nx5271, CLK=>clk, 
      R=>nx14156);
   booth_integrtaion_5_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_5, QB=>OPEN, D=>nx5261, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_5, QB=>OPEN, D=>nx5251, CLK=>clk, 
      R=>nx14154);
   booth_integrtaion_5_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_4, QB=>OPEN, D=>nx5241, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_4, QB=>OPEN, D=>nx5231, CLK=>clk, 
      R=>nx14154);
   booth_integrtaion_5_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_3, QB=>OPEN, D=>nx5221, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_3, QB=>OPEN, D=>nx5211, CLK=>clk, 
      R=>nx14154);
   booth_integrtaion_5_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_2, QB=>OPEN, D=>nx5201, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_2, QB=>OPEN, D=>nx5191, CLK=>clk, 
      R=>nx14154);
   booth_integrtaion_5_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_output_1, QB=>OPEN, D=>nx5181, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_5_shift_Reg_count_1, QB=>OPEN, D=>nx5171, CLK=>clk, 
      R=>nx14154);
   ix5142 : nand02 port map ( Y=>nx5141, A0=>nx14628, A1=>nx14248);
   booth_integrtaion_5_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx11075, D=>nx5141, CLK=>clk, S=>nx14154);
   ix4587 : nand02 port map ( Y=>nx4586, A0=>nx11096, A1=>nx11107);
   ix11097 : oai21 port map ( Y=>nx11096, A0=>nx4050, A1=>nx4046, B0=>
      weight_5(0));
   ix5352 : oai21 port map ( Y=>nx5351, A0=>nx11101, A1=>nx14476, B0=>
      nx11103);
   booth_integrtaion_5_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11101, D=>nx5351, CLK=>clk, R=>rst);
   booth_integrtaion_5_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_0, QB=>nx10980, D=>nx5661, CLK=>clk, R=>rst
   );
   ix11112 : xnor2 port map ( Y=>nx11111, A0=>nx4056, A1=>nx2921);
   ix5492 : oai21 port map ( Y=>nx5491, A0=>nx11117, A1=>nx14476, B0=>
      nx11119);
   booth_integrtaion_5_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_17, QB=>nx11117, D=>nx5491, CLK=>clk, 
      R=>rst);
   ix11120 : nand03 port map ( Y=>nx11119, A0=>nx14484, A1=>nx4564, A2=>
      nx14722);
   ix4565 : xnor2 port map ( Y=>nx4564, A0=>nx11122, A1=>nx2923);
   ix11123 : aoi22 port map ( Y=>nx11122, A0=>
      booth_integrtaion_5_booth_output_17, A1=>nx4080, B0=>nx4056, B1=>
      nx2921);
   ix4065 : nand02 port map ( Y=>nx4064, A0=>weight_5(1), A1=>weight_5(0));
   ix11127 : or02 port map ( Y=>nx11126, A0=>weight_5(0), A1=>weight_5(1));
   ix5482 : oai21 port map ( Y=>nx5481, A0=>nx11131, A1=>nx14476, B0=>
      nx11133);
   booth_integrtaion_5_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11131, D=>nx5481, CLK=>clk, R=>rst);
   ix11134 : nand03 port map ( Y=>nx11133, A0=>nx14484, A1=>nx4552, A2=>
      nx14722);
   ix4553 : xnor2 port map ( Y=>nx4552, A0=>nx4108, A1=>nx11144);
   ix4109 : oai22 port map ( Y=>nx4108, A0=>nx11122, A1=>nx11137, B0=>
      nx11131, B1=>nx14488);
   ix11140 : aoi32 port map ( Y=>nx11139, A0=>nx4090, A1=>nx4050, A2=>
      nx11142, B0=>weight_5(2), B1=>nx4046);
   ix4091 : oai21 port map ( Y=>nx4090, A0=>weight_5(0), A1=>weight_5(1), B0
      =>weight_5(2));
   ix11145 : xnor2 port map ( Y=>nx11144, A0=>
      booth_integrtaion_5_booth_output_19, A1=>nx4128);
   booth_integrtaion_5_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_19, QB=>OPEN, D=>nx5471, CLK=>clk, R
      =>rst);
   ix11150 : xnor2 port map ( Y=>nx11149, A0=>nx11151, A1=>nx11165);
   ix11152 : aoi22 port map ( Y=>nx11151, A0=>
      booth_integrtaion_5_booth_output_19, A1=>nx4128, B0=>nx4108, B1=>
      nx2925);
   ix4129 : oai32 port map ( Y=>nx4128, A0=>nx11154, A1=>nx14490, A2=>nx4118, 
      B0=>nx11160, B1=>nx14494);
   ix11155 : nor02ii port map ( Y=>nx11154, A0=>nx4094, A1=>weight_5(3));
   ix4095 : nor03_2x port map ( Y=>nx4094, A0=>weight_5(2), A1=>weight_5(0), 
      A2=>weight_5(1));
   ix4119 : nor04 port map ( Y=>nx4118, A0=>weight_5(3), A1=>weight_5(2), A2
      =>weight_5(0), A3=>weight_5(1));
   ix11161 : inv01 port map ( Y=>nx11160, A=>weight_5(3));
   ix5462 : oai21 port map ( Y=>nx5461, A0=>nx11169, A1=>nx14476, B0=>
      nx11171);
   booth_integrtaion_5_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11169, D=>nx5461, CLK=>clk, R=>rst);
   ix11172 : nand03 port map ( Y=>nx11171, A0=>nx14484, A1=>nx4528, A2=>
      nx14722);
   ix4529 : xnor2 port map ( Y=>nx4528, A0=>nx4156, A1=>nx11184);
   ix4157 : oai22 port map ( Y=>nx4156, A0=>nx11151, A1=>nx11165, B0=>
      nx11169, B1=>nx11175);
   ix11183 : inv01 port map ( Y=>nx11182, A=>weight_5(4));
   ix11185 : xnor2 port map ( Y=>nx11184, A0=>
      booth_integrtaion_5_booth_output_21, A1=>nx4176);
   booth_integrtaion_5_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_21, QB=>OPEN, D=>nx5451, CLK=>clk, R
      =>rst);
   ix11190 : xnor2 port map ( Y=>nx11189, A0=>nx11191, A1=>nx11201);
   ix11192 : aoi22 port map ( Y=>nx11191, A0=>
      booth_integrtaion_5_booth_output_21, A1=>nx4176, B0=>nx4156, B1=>
      nx2928);
   ix4177 : oai32 port map ( Y=>nx4176, A0=>nx11194, A1=>nx14490, A2=>nx4166, 
      B0=>nx11198, B1=>nx14494);
   ix11195 : nor02ii port map ( Y=>nx11194, A0=>nx4142, A1=>weight_5(5));
   ix4143 : nor02ii port map ( Y=>nx4142, A0=>weight_5(4), A1=>nx4118);
   ix4167 : nor02ii port map ( Y=>nx4166, A0=>weight_5(5), A1=>nx4142);
   ix11199 : inv01 port map ( Y=>nx11198, A=>weight_5(5));
   ix5442 : oai21 port map ( Y=>nx5441, A0=>nx11205, A1=>nx14476, B0=>
      nx11207);
   booth_integrtaion_5_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11205, D=>nx5441, CLK=>clk, R=>rst);
   ix11208 : nand03 port map ( Y=>nx11207, A0=>nx14484, A1=>nx4504, A2=>
      nx14478);
   ix4505 : xnor2 port map ( Y=>nx4504, A0=>nx4204, A1=>nx11220);
   ix4205 : oai22 port map ( Y=>nx4204, A0=>nx11191, A1=>nx11201, B0=>
      nx11205, B1=>nx11211);
   ix11219 : inv01 port map ( Y=>nx11218, A=>weight_5(6));
   ix11221 : xnor2 port map ( Y=>nx11220, A0=>
      booth_integrtaion_5_booth_output_23, A1=>nx4224);
   booth_integrtaion_5_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_23, QB=>OPEN, D=>nx5431, CLK=>clk, R
      =>rst);
   ix11226 : xnor2 port map ( Y=>nx11225, A0=>nx11227, A1=>nx11237);
   ix11228 : aoi22 port map ( Y=>nx11227, A0=>
      booth_integrtaion_5_booth_output_23, A1=>nx4224, B0=>nx4204, B1=>
      nx2930);
   ix4225 : oai32 port map ( Y=>nx4224, A0=>nx11230, A1=>nx14490, A2=>nx4214, 
      B0=>nx11234, B1=>nx14494);
   ix11231 : nor02ii port map ( Y=>nx11230, A0=>nx4190, A1=>weight_5(7));
   ix4191 : nor02ii port map ( Y=>nx4190, A0=>weight_5(6), A1=>nx4166);
   ix4215 : nor02ii port map ( Y=>nx4214, A0=>weight_5(7), A1=>nx4190);
   ix11235 : inv01 port map ( Y=>nx11234, A=>weight_5(7));
   ix5422 : oai21 port map ( Y=>nx5421, A0=>nx11241, A1=>nx14478, B0=>
      nx11243);
   booth_integrtaion_5_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11241, D=>nx5421, CLK=>clk, R=>rst);
   ix11244 : nand03 port map ( Y=>nx11243, A0=>nx14484, A1=>nx4480, A2=>
      nx14478);
   ix4481 : xnor2 port map ( Y=>nx4480, A0=>nx4252, A1=>nx11256);
   ix4253 : oai22 port map ( Y=>nx4252, A0=>nx11227, A1=>nx11237, B0=>
      nx11241, B1=>nx11247);
   ix11255 : inv01 port map ( Y=>nx11254, A=>weight_5(8));
   ix11257 : xnor2 port map ( Y=>nx11256, A0=>
      booth_integrtaion_5_booth_output_25, A1=>nx4272);
   booth_integrtaion_5_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_25, QB=>OPEN, D=>nx5411, CLK=>clk, R
      =>rst);
   ix11262 : xnor2 port map ( Y=>nx11261, A0=>nx11263, A1=>nx11273);
   ix11264 : aoi22 port map ( Y=>nx11263, A0=>
      booth_integrtaion_5_booth_output_25, A1=>nx4272, B0=>nx4252, B1=>
      nx2932);
   ix4273 : oai32 port map ( Y=>nx4272, A0=>nx11266, A1=>nx14490, A2=>nx4262, 
      B0=>nx11270, B1=>nx14494);
   ix11267 : nor02ii port map ( Y=>nx11266, A0=>nx4238, A1=>weight_5(9));
   ix4239 : nor02ii port map ( Y=>nx4238, A0=>weight_5(8), A1=>nx4214);
   ix4263 : nor02ii port map ( Y=>nx4262, A0=>weight_5(9), A1=>nx4238);
   ix11271 : inv01 port map ( Y=>nx11270, A=>weight_5(9));
   ix5402 : oai21 port map ( Y=>nx5401, A0=>nx11277, A1=>nx14478, B0=>
      nx11279);
   booth_integrtaion_5_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11277, D=>nx5401, CLK=>clk, R=>rst);
   ix11280 : nand03 port map ( Y=>nx11279, A0=>nx14484, A1=>nx4456, A2=>
      nx14478);
   ix4457 : xnor2 port map ( Y=>nx4456, A0=>nx4300, A1=>nx11292);
   ix4301 : oai22 port map ( Y=>nx4300, A0=>nx11263, A1=>nx11273, B0=>
      nx11277, B1=>nx11283);
   ix11291 : inv01 port map ( Y=>nx11290, A=>weight_5(10));
   ix11293 : xnor2 port map ( Y=>nx11292, A0=>
      booth_integrtaion_5_booth_output_27, A1=>nx4320);
   booth_integrtaion_5_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_27, QB=>OPEN, D=>nx5391, CLK=>clk, R
      =>rst);
   ix11298 : xnor2 port map ( Y=>nx11297, A0=>nx11299, A1=>nx11309);
   ix11300 : aoi22 port map ( Y=>nx11299, A0=>
      booth_integrtaion_5_booth_output_27, A1=>nx4320, B0=>nx4300, B1=>
      nx2934);
   ix4321 : oai32 port map ( Y=>nx4320, A0=>nx11302, A1=>nx14490, A2=>nx4310, 
      B0=>nx11306, B1=>nx14494);
   ix11303 : nor02ii port map ( Y=>nx11302, A0=>nx4286, A1=>weight_5(11));
   ix4287 : nor02ii port map ( Y=>nx4286, A0=>weight_5(10), A1=>nx4262);
   ix4311 : nor02ii port map ( Y=>nx4310, A0=>weight_5(11), A1=>nx4286);
   ix11307 : inv01 port map ( Y=>nx11306, A=>weight_5(11));
   ix5382 : oai21 port map ( Y=>nx5381, A0=>nx11313, A1=>nx14478, B0=>
      nx11315);
   booth_integrtaion_5_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11313, D=>nx5381, CLK=>clk, R=>rst);
   ix11316 : nand03 port map ( Y=>nx11315, A0=>nx14730, A1=>nx4432, A2=>
      nx14478);
   ix4433 : xnor2 port map ( Y=>nx4432, A0=>nx4348, A1=>nx11328);
   ix4349 : oai22 port map ( Y=>nx4348, A0=>nx11299, A1=>nx11309, B0=>
      nx11313, B1=>nx11319);
   ix11327 : inv01 port map ( Y=>nx11326, A=>weight_5(12));
   ix11329 : xnor2 port map ( Y=>nx11328, A0=>
      booth_integrtaion_5_booth_output_29, A1=>nx4368);
   booth_integrtaion_5_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_29, QB=>OPEN, D=>nx5371, CLK=>clk, R
      =>rst);
   ix11334 : xnor2 port map ( Y=>nx11333, A0=>nx11335, A1=>nx11345);
   ix11336 : aoi22 port map ( Y=>nx11335, A0=>
      booth_integrtaion_5_booth_output_29, A1=>nx4368, B0=>nx4348, B1=>
      nx2936);
   ix4369 : oai32 port map ( Y=>nx4368, A0=>nx11338, A1=>nx14490, A2=>nx4358, 
      B0=>nx11342, B1=>nx14494);
   ix11339 : nor02ii port map ( Y=>nx11338, A0=>nx4334, A1=>weight_5(13));
   ix4335 : nor02ii port map ( Y=>nx4334, A0=>weight_5(12), A1=>nx4310);
   ix4359 : nor02ii port map ( Y=>nx4358, A0=>weight_5(13), A1=>nx4334);
   ix11343 : inv01 port map ( Y=>nx11342, A=>weight_5(13));
   ix11351 : xnor2 port map ( Y=>nx11350, A0=>nx4396, A1=>nx4406);
   ix4397 : oai22 port map ( Y=>nx4396, A0=>nx11335, A1=>nx11345, B0=>
      nx11353, B1=>nx11355);
   booth_integrtaion_5_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_31, QB=>nx11353, D=>nx5361, CLK=>clk, 
      R=>rst);
   ix11363 : inv01 port map ( Y=>nx11362, A=>weight_5(14));
   ix11366 : aoi22 port map ( Y=>nx11365, A0=>weight_5(15), A1=>nx4046, B0=>
      nx4050, B1=>nx4398);
   ix4399 : xnor2 port map ( Y=>nx4398, A0=>weight_5(15), A1=>nx4382);
   ix4383 : nor02ii port map ( Y=>nx4382, A0=>weight_5(14), A1=>nx4358);
   ix4393 : oai32 port map ( Y=>nx4392, A0=>nx11370, A1=>nx14490, A2=>nx4382, 
      B0=>nx11362, B1=>nx14494);
   ix11371 : nor02ii port map ( Y=>nx11370, A0=>nx4358, A1=>weight_5(14));
   ix4345 : oai32 port map ( Y=>nx4344, A0=>nx11374, A1=>nx14492, A2=>nx4334, 
      B0=>nx11326, B1=>nx14496);
   ix11375 : nor02ii port map ( Y=>nx11374, A0=>nx4310, A1=>weight_5(12));
   ix4297 : oai32 port map ( Y=>nx4296, A0=>nx11378, A1=>nx14492, A2=>nx4286, 
      B0=>nx11290, B1=>nx14496);
   ix11379 : nor02ii port map ( Y=>nx11378, A0=>nx4262, A1=>weight_5(10));
   ix4249 : oai32 port map ( Y=>nx4248, A0=>nx11382, A1=>nx14492, A2=>nx4238, 
      B0=>nx11254, B1=>nx14496);
   ix11383 : nor02ii port map ( Y=>nx11382, A0=>nx4214, A1=>weight_5(8));
   ix4201 : oai32 port map ( Y=>nx4200, A0=>nx11386, A1=>nx14492, A2=>nx4190, 
      B0=>nx11218, B1=>nx14496);
   ix11387 : nor02ii port map ( Y=>nx11386, A0=>nx4166, A1=>weight_5(6));
   ix4153 : oai32 port map ( Y=>nx4152, A0=>nx11390, A1=>nx14492, A2=>nx4142, 
      B0=>nx11182, B1=>nx14496);
   ix11391 : nor02ii port map ( Y=>nx11390, A0=>nx4118, A1=>weight_5(4));
   ix11394 : aoi32 port map ( Y=>nx11393, A0=>nx4064, A1=>nx4050, A2=>
      nx11126, B0=>weight_5(1), B1=>nx4046);
   booth_integrtaion_5_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_5_booth_output_16, QB=>nx11107, D=>nx5501, CLK=>clk, 
      R=>rst);
   booth_integrtaion_5_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_5_15, QB=>nx11397, D=>nx5511, CLK=>clk, R=>
      rst);
   ix4929 : xor2 port map ( Y=>label_5(1), A0=>nx11414, A1=>nx11416);
   ix11415 : nand02 port map ( Y=>nx11414, A0=>adderInput_5(0), A1=>
      booth_integration_output_5_0);
   ix11417 : xnor2 port map ( Y=>nx11416, A0=>booth_integration_output_5_1, 
      A1=>adderInput_5(1));
   ix4927 : xor2 port map ( Y=>label_5(2), A0=>nx11419, A1=>nx11422);
   ix11420 : aoi32 port map ( Y=>nx11419, A0=>adderInput_5(0), A1=>
      booth_integration_output_5_0, A2=>nx4786, B0=>adderInput_5(1), B1=>
      booth_integration_output_5_1);
   ix4925 : xnor2 port map ( Y=>label_5(3), A0=>nx4800, A1=>nx11428);
   ix4801 : oai22 port map ( Y=>nx4800, A0=>nx11419, A1=>nx11422, B0=>
      nx11426, B1=>nx11411);
   ix11427 : inv01 port map ( Y=>nx11426, A=>adderInput_5(2));
   ix11429 : xnor2 port map ( Y=>nx11428, A0=>booth_integration_output_5_3, 
      A1=>adderInput_5(3));
   ix4923 : xor2 port map ( Y=>label_5(4), A0=>nx11431, A1=>nx11434);
   ix11432 : aoi22 port map ( Y=>nx11431, A0=>adderInput_5(3), A1=>
      booth_integration_output_5_3, B0=>nx4800, B1=>nx4802);
   ix4921 : xnor2 port map ( Y=>label_5(5), A0=>nx4816, A1=>nx11440);
   ix4817 : oai22 port map ( Y=>nx4816, A0=>nx11431, A1=>nx11434, B0=>
      nx11438, B1=>nx11409);
   ix11439 : inv01 port map ( Y=>nx11438, A=>adderInput_5(4));
   ix11441 : xnor2 port map ( Y=>nx11440, A0=>booth_integration_output_5_5, 
      A1=>adderInput_5(5));
   ix4919 : xor2 port map ( Y=>label_5(6), A0=>nx11443, A1=>nx11446);
   ix11444 : aoi22 port map ( Y=>nx11443, A0=>adderInput_5(5), A1=>
      booth_integration_output_5_5, B0=>nx4816, B1=>nx4818);
   ix4917 : xnor2 port map ( Y=>label_5(7), A0=>nx4832, A1=>nx11452);
   ix4833 : oai22 port map ( Y=>nx4832, A0=>nx11443, A1=>nx11446, B0=>
      nx11450, B1=>nx11407);
   ix11451 : inv01 port map ( Y=>nx11450, A=>adderInput_5(6));
   ix11453 : xnor2 port map ( Y=>nx11452, A0=>booth_integration_output_5_7, 
      A1=>adderInput_5(7));
   ix4915 : xor2 port map ( Y=>label_5(8), A0=>nx11455, A1=>nx11458);
   ix11456 : aoi22 port map ( Y=>nx11455, A0=>adderInput_5(7), A1=>
      booth_integration_output_5_7, B0=>nx4832, B1=>nx4834);
   ix4913 : xnor2 port map ( Y=>label_5(9), A0=>nx4848, A1=>nx11464);
   ix4849 : oai22 port map ( Y=>nx4848, A0=>nx11455, A1=>nx11458, B0=>
      nx11462, B1=>nx11405);
   ix11463 : inv01 port map ( Y=>nx11462, A=>adderInput_5(8));
   ix11465 : xnor2 port map ( Y=>nx11464, A0=>booth_integration_output_5_9, 
      A1=>adderInput_5(9));
   ix4911 : xor2 port map ( Y=>label_5(10), A0=>nx11467, A1=>nx11470);
   ix11468 : aoi22 port map ( Y=>nx11467, A0=>adderInput_5(9), A1=>
      booth_integration_output_5_9, B0=>nx4848, B1=>nx4850);
   ix4909 : xnor2 port map ( Y=>label_5(11), A0=>nx4864, A1=>nx11476);
   ix4865 : oai22 port map ( Y=>nx4864, A0=>nx11467, A1=>nx11470, B0=>
      nx11474, B1=>nx11403);
   ix11475 : inv01 port map ( Y=>nx11474, A=>adderInput_5(10));
   ix11477 : xnor2 port map ( Y=>nx11476, A0=>booth_integration_output_5_11, 
      A1=>adderInput_5(11));
   ix4907 : xor2 port map ( Y=>label_5(12), A0=>nx11479, A1=>nx11482);
   ix11480 : aoi22 port map ( Y=>nx11479, A0=>adderInput_5(11), A1=>
      booth_integration_output_5_11, B0=>nx4864, B1=>nx4866);
   ix4905 : xnor2 port map ( Y=>label_5(13), A0=>nx4880, A1=>nx11488);
   ix4881 : oai22 port map ( Y=>nx4880, A0=>nx11479, A1=>nx11482, B0=>
      nx11486, B1=>nx11401);
   ix11487 : inv01 port map ( Y=>nx11486, A=>adderInput_5(12));
   ix11489 : xnor2 port map ( Y=>nx11488, A0=>booth_integration_output_5_13, 
      A1=>adderInput_5(13));
   ix4903 : xor2 port map ( Y=>label_5(14), A0=>nx11491, A1=>nx11494);
   ix11492 : aoi22 port map ( Y=>nx11491, A0=>adderInput_5(13), A1=>
      booth_integration_output_5_13, B0=>nx4880, B1=>nx4882);
   ix4901 : xnor2 port map ( Y=>label_5(15), A0=>nx4896, A1=>nx11500);
   ix4897 : oai22 port map ( Y=>nx4896, A0=>nx11491, A1=>nx11494, B0=>
      nx11498, B1=>nx11399);
   ix11499 : inv01 port map ( Y=>nx11498, A=>adderInput_5(14));
   booth_integrtaion_4_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_1, QB=>OPEN, D=>nx6181, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_2, QB=>nx11934, D=>nx6171, CLK=>clk, R=>rst
   );
   booth_integrtaion_4_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_3, QB=>OPEN, D=>nx6161, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_4, QB=>nx11932, D=>nx6151, CLK=>clk, R=>rst
   );
   booth_integrtaion_4_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_5, QB=>OPEN, D=>nx6141, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_6, QB=>nx11930, D=>nx6131, CLK=>clk, R=>rst
   );
   booth_integrtaion_4_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_7, QB=>OPEN, D=>nx6121, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_8, QB=>nx11928, D=>nx6111, CLK=>clk, R=>rst
   );
   booth_integrtaion_4_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_9, QB=>OPEN, D=>nx6101, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_10, QB=>nx11926, D=>nx6091, CLK=>clk, R=>
      rst);
   booth_integrtaion_4_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_11, QB=>OPEN, D=>nx6081, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_12, QB=>nx11924, D=>nx6071, CLK=>clk, R=>
      rst);
   booth_integrtaion_4_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_13, QB=>OPEN, D=>nx6061, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_14, QB=>nx11922, D=>nx6051, CLK=>clk, R=>
      rst);
   ix11552 : aoi22 port map ( Y=>nx11551, A0=>neuron(15), A1=>nx14284, B0=>
      nx5572, B1=>nx5578);
   booth_integrtaion_4_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_reg_output_0, QB=>OPEN, D=>nx5691, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_0, QB=>OPEN, D=>nx5677, CLK=>clk, 
      S=>nx14160);
   booth_integrtaion_4_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_reg_output_9, QB=>OPEN, D=>nx5871, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_9, QB=>OPEN, D=>nx5861, CLK=>clk, 
      R=>nx14160);
   booth_integrtaion_4_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_8, QB=>OPEN, D=>nx5851, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_8, QB=>OPEN, D=>nx5841, CLK=>clk, 
      R=>nx14158);
   booth_integrtaion_4_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_7, QB=>OPEN, D=>nx5831, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_7, QB=>OPEN, D=>nx5821, CLK=>clk, 
      R=>nx14158);
   booth_integrtaion_4_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_6, QB=>OPEN, D=>nx5811, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_6, QB=>OPEN, D=>nx5801, CLK=>clk, 
      R=>nx14158);
   booth_integrtaion_4_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_5, QB=>OPEN, D=>nx5791, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_5, QB=>OPEN, D=>nx5781, CLK=>clk, 
      R=>nx14158);
   booth_integrtaion_4_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_4, QB=>OPEN, D=>nx5771, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_4, QB=>OPEN, D=>nx5761, CLK=>clk, 
      R=>nx14158);
   booth_integrtaion_4_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_3, QB=>OPEN, D=>nx5751, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_3, QB=>OPEN, D=>nx5741, CLK=>clk, 
      R=>nx14158);
   booth_integrtaion_4_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_2, QB=>OPEN, D=>nx5731, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_2, QB=>OPEN, D=>nx5721, CLK=>clk, 
      R=>nx14158);
   booth_integrtaion_4_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_output_1, QB=>OPEN, D=>nx5711, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_4_shift_Reg_count_1, QB=>OPEN, D=>nx5701, CLK=>clk, 
      R=>nx14156);
   ix5672 : nand02 port map ( Y=>nx5671, A0=>nx14632, A1=>nx14270);
   booth_integrtaion_4_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx11598, D=>nx5671, CLK=>clk, S=>nx14156);
   ix5573 : nand02 port map ( Y=>nx5572, A0=>nx11619, A1=>nx11630);
   ix11620 : oai21 port map ( Y=>nx11619, A0=>nx5036, A1=>nx5032, B0=>
      weight_4(0));
   ix5882 : oai21 port map ( Y=>nx5881, A0=>nx11624, A1=>nx14498, B0=>
      nx11626);
   booth_integrtaion_4_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11624, D=>nx5881, CLK=>clk, R=>rst);
   booth_integrtaion_4_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_0, QB=>nx11503, D=>nx6191, CLK=>clk, R=>rst
   );
   ix11635 : xnor2 port map ( Y=>nx11634, A0=>nx5042, A1=>nx2939);
   ix6022 : oai21 port map ( Y=>nx6021, A0=>nx11640, A1=>nx14498, B0=>
      nx11642);
   booth_integrtaion_4_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_17, QB=>nx11640, D=>nx6021, CLK=>clk, 
      R=>rst);
   ix11643 : nand03 port map ( Y=>nx11642, A0=>nx14506, A1=>nx5550, A2=>
      nx14738);
   ix5551 : xnor2 port map ( Y=>nx5550, A0=>nx11645, A1=>nx2940);
   ix11646 : aoi22 port map ( Y=>nx11645, A0=>
      booth_integrtaion_4_booth_output_17, A1=>nx5066, B0=>nx5042, B1=>
      nx2939);
   ix5051 : nand02 port map ( Y=>nx5050, A0=>weight_4(1), A1=>weight_4(0));
   ix11650 : or02 port map ( Y=>nx11649, A0=>weight_4(0), A1=>weight_4(1));
   ix6012 : oai21 port map ( Y=>nx6011, A0=>nx11654, A1=>nx14498, B0=>
      nx11656);
   booth_integrtaion_4_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11654, D=>nx6011, CLK=>clk, R=>rst);
   ix11657 : nand03 port map ( Y=>nx11656, A0=>nx14506, A1=>nx5538, A2=>
      nx14738);
   ix5539 : xnor2 port map ( Y=>nx5538, A0=>nx5094, A1=>nx11667);
   ix5095 : oai22 port map ( Y=>nx5094, A0=>nx11645, A1=>nx11660, B0=>
      nx11654, B1=>nx14510);
   ix11663 : aoi32 port map ( Y=>nx11662, A0=>nx5076, A1=>nx5036, A2=>
      nx11665, B0=>weight_4(2), B1=>nx5032);
   ix5077 : oai21 port map ( Y=>nx5076, A0=>weight_4(0), A1=>weight_4(1), B0
      =>weight_4(2));
   ix11668 : xnor2 port map ( Y=>nx11667, A0=>
      booth_integrtaion_4_booth_output_19, A1=>nx5114);
   booth_integrtaion_4_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_19, QB=>OPEN, D=>nx6001, CLK=>clk, R
      =>rst);
   ix11673 : xnor2 port map ( Y=>nx11672, A0=>nx11674, A1=>nx11688);
   ix11675 : aoi22 port map ( Y=>nx11674, A0=>
      booth_integrtaion_4_booth_output_19, A1=>nx5114, B0=>nx5094, B1=>
      nx2941);
   ix5115 : oai32 port map ( Y=>nx5114, A0=>nx11677, A1=>nx14512, A2=>nx5104, 
      B0=>nx11683, B1=>nx14516);
   ix11678 : nor02ii port map ( Y=>nx11677, A0=>nx5080, A1=>weight_4(3));
   ix5081 : nor03_2x port map ( Y=>nx5080, A0=>weight_4(2), A1=>weight_4(0), 
      A2=>weight_4(1));
   ix5105 : nor04 port map ( Y=>nx5104, A0=>weight_4(3), A1=>weight_4(2), A2
      =>weight_4(0), A3=>weight_4(1));
   ix11684 : inv01 port map ( Y=>nx11683, A=>weight_4(3));
   ix5992 : oai21 port map ( Y=>nx5991, A0=>nx11692, A1=>nx14498, B0=>
      nx11694);
   booth_integrtaion_4_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11692, D=>nx5991, CLK=>clk, R=>rst);
   ix11695 : nand03 port map ( Y=>nx11694, A0=>nx14506, A1=>nx5514, A2=>
      nx14738);
   ix5515 : xnor2 port map ( Y=>nx5514, A0=>nx5142, A1=>nx11707);
   ix5143 : oai22 port map ( Y=>nx5142, A0=>nx11674, A1=>nx11688, B0=>
      nx11692, B1=>nx11698);
   ix11706 : inv01 port map ( Y=>nx11705, A=>weight_4(4));
   ix11708 : xnor2 port map ( Y=>nx11707, A0=>
      booth_integrtaion_4_booth_output_21, A1=>nx5162);
   booth_integrtaion_4_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_21, QB=>OPEN, D=>nx5981, CLK=>clk, R
      =>rst);
   ix11713 : xnor2 port map ( Y=>nx11712, A0=>nx11714, A1=>nx11724);
   ix11715 : aoi22 port map ( Y=>nx11714, A0=>
      booth_integrtaion_4_booth_output_21, A1=>nx5162, B0=>nx5142, B1=>
      nx2943);
   ix5163 : oai32 port map ( Y=>nx5162, A0=>nx11717, A1=>nx14512, A2=>nx5152, 
      B0=>nx11721, B1=>nx14516);
   ix11718 : nor02ii port map ( Y=>nx11717, A0=>nx5128, A1=>weight_4(5));
   ix5129 : nor02ii port map ( Y=>nx5128, A0=>weight_4(4), A1=>nx5104);
   ix5153 : nor02ii port map ( Y=>nx5152, A0=>weight_4(5), A1=>nx5128);
   ix11722 : inv01 port map ( Y=>nx11721, A=>weight_4(5));
   ix5972 : oai21 port map ( Y=>nx5971, A0=>nx11728, A1=>nx14498, B0=>
      nx11730);
   booth_integrtaion_4_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11728, D=>nx5971, CLK=>clk, R=>rst);
   ix11731 : nand03 port map ( Y=>nx11730, A0=>nx14506, A1=>nx5490, A2=>
      nx14500);
   ix5491 : xnor2 port map ( Y=>nx5490, A0=>nx5190, A1=>nx11743);
   ix5191 : oai22 port map ( Y=>nx5190, A0=>nx11714, A1=>nx11724, B0=>
      nx11728, B1=>nx11734);
   ix11742 : inv01 port map ( Y=>nx11741, A=>weight_4(6));
   ix11744 : xnor2 port map ( Y=>nx11743, A0=>
      booth_integrtaion_4_booth_output_23, A1=>nx5210);
   booth_integrtaion_4_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_23, QB=>OPEN, D=>nx5961, CLK=>clk, R
      =>rst);
   ix11749 : xnor2 port map ( Y=>nx11748, A0=>nx11750, A1=>nx11760);
   ix11751 : aoi22 port map ( Y=>nx11750, A0=>
      booth_integrtaion_4_booth_output_23, A1=>nx5210, B0=>nx5190, B1=>
      nx2945);
   ix5211 : oai32 port map ( Y=>nx5210, A0=>nx11753, A1=>nx14512, A2=>nx5200, 
      B0=>nx11757, B1=>nx14516);
   ix11754 : nor02ii port map ( Y=>nx11753, A0=>nx5176, A1=>weight_4(7));
   ix5177 : nor02ii port map ( Y=>nx5176, A0=>weight_4(6), A1=>nx5152);
   ix5201 : nor02ii port map ( Y=>nx5200, A0=>weight_4(7), A1=>nx5176);
   ix11758 : inv01 port map ( Y=>nx11757, A=>weight_4(7));
   ix5952 : oai21 port map ( Y=>nx5951, A0=>nx11764, A1=>nx14500, B0=>
      nx11766);
   booth_integrtaion_4_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11764, D=>nx5951, CLK=>clk, R=>rst);
   ix11767 : nand03 port map ( Y=>nx11766, A0=>nx14506, A1=>nx5466, A2=>
      nx14500);
   ix5467 : xnor2 port map ( Y=>nx5466, A0=>nx5238, A1=>nx11779);
   ix5239 : oai22 port map ( Y=>nx5238, A0=>nx11750, A1=>nx11760, B0=>
      nx11764, B1=>nx11770);
   ix11778 : inv01 port map ( Y=>nx11777, A=>weight_4(8));
   ix11780 : xnor2 port map ( Y=>nx11779, A0=>
      booth_integrtaion_4_booth_output_25, A1=>nx5258);
   booth_integrtaion_4_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_25, QB=>OPEN, D=>nx5941, CLK=>clk, R
      =>rst);
   ix11785 : xnor2 port map ( Y=>nx11784, A0=>nx11786, A1=>nx11796);
   ix11787 : aoi22 port map ( Y=>nx11786, A0=>
      booth_integrtaion_4_booth_output_25, A1=>nx5258, B0=>nx5238, B1=>
      nx2947);
   ix5259 : oai32 port map ( Y=>nx5258, A0=>nx11789, A1=>nx14512, A2=>nx5248, 
      B0=>nx11793, B1=>nx14516);
   ix11790 : nor02ii port map ( Y=>nx11789, A0=>nx5224, A1=>weight_4(9));
   ix5225 : nor02ii port map ( Y=>nx5224, A0=>weight_4(8), A1=>nx5200);
   ix5249 : nor02ii port map ( Y=>nx5248, A0=>weight_4(9), A1=>nx5224);
   ix11794 : inv01 port map ( Y=>nx11793, A=>weight_4(9));
   ix5932 : oai21 port map ( Y=>nx5931, A0=>nx11800, A1=>nx14500, B0=>
      nx11802);
   booth_integrtaion_4_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11800, D=>nx5931, CLK=>clk, R=>rst);
   ix11803 : nand03 port map ( Y=>nx11802, A0=>nx14506, A1=>nx5442, A2=>
      nx14500);
   ix5443 : xnor2 port map ( Y=>nx5442, A0=>nx5286, A1=>nx11815);
   ix5287 : oai22 port map ( Y=>nx5286, A0=>nx11786, A1=>nx11796, B0=>
      nx11800, B1=>nx11806);
   ix11814 : inv01 port map ( Y=>nx11813, A=>weight_4(10));
   ix11816 : xnor2 port map ( Y=>nx11815, A0=>
      booth_integrtaion_4_booth_output_27, A1=>nx5306);
   booth_integrtaion_4_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_27, QB=>OPEN, D=>nx5921, CLK=>clk, R
      =>rst);
   ix11821 : xnor2 port map ( Y=>nx11820, A0=>nx11822, A1=>nx11832);
   ix11823 : aoi22 port map ( Y=>nx11822, A0=>
      booth_integrtaion_4_booth_output_27, A1=>nx5306, B0=>nx5286, B1=>
      nx2949);
   ix5307 : oai32 port map ( Y=>nx5306, A0=>nx11825, A1=>nx14512, A2=>nx5296, 
      B0=>nx11829, B1=>nx14516);
   ix11826 : nor02ii port map ( Y=>nx11825, A0=>nx5272, A1=>weight_4(11));
   ix5273 : nor02ii port map ( Y=>nx5272, A0=>weight_4(10), A1=>nx5248);
   ix5297 : nor02ii port map ( Y=>nx5296, A0=>weight_4(11), A1=>nx5272);
   ix11830 : inv01 port map ( Y=>nx11829, A=>weight_4(11));
   ix5912 : oai21 port map ( Y=>nx5911, A0=>nx11836, A1=>nx14500, B0=>
      nx11838);
   booth_integrtaion_4_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx11836, D=>nx5911, CLK=>clk, R=>rst);
   ix11839 : nand03 port map ( Y=>nx11838, A0=>nx14746, A1=>nx5418, A2=>
      nx14500);
   ix5419 : xnor2 port map ( Y=>nx5418, A0=>nx5334, A1=>nx11851);
   ix5335 : oai22 port map ( Y=>nx5334, A0=>nx11822, A1=>nx11832, B0=>
      nx11836, B1=>nx11842);
   ix11850 : inv01 port map ( Y=>nx11849, A=>weight_4(12));
   ix11852 : xnor2 port map ( Y=>nx11851, A0=>
      booth_integrtaion_4_booth_output_29, A1=>nx5354);
   booth_integrtaion_4_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_29, QB=>OPEN, D=>nx5901, CLK=>clk, R
      =>rst);
   ix11857 : xnor2 port map ( Y=>nx11856, A0=>nx11858, A1=>nx11868);
   ix11859 : aoi22 port map ( Y=>nx11858, A0=>
      booth_integrtaion_4_booth_output_29, A1=>nx5354, B0=>nx5334, B1=>
      nx2951);
   ix5355 : oai32 port map ( Y=>nx5354, A0=>nx11861, A1=>nx14512, A2=>nx5344, 
      B0=>nx11865, B1=>nx14516);
   ix11862 : nor02ii port map ( Y=>nx11861, A0=>nx5320, A1=>weight_4(13));
   ix5321 : nor02ii port map ( Y=>nx5320, A0=>weight_4(12), A1=>nx5296);
   ix5345 : nor02ii port map ( Y=>nx5344, A0=>weight_4(13), A1=>nx5320);
   ix11866 : inv01 port map ( Y=>nx11865, A=>weight_4(13));
   ix11874 : xnor2 port map ( Y=>nx11873, A0=>nx5382, A1=>nx5392);
   ix5383 : oai22 port map ( Y=>nx5382, A0=>nx11858, A1=>nx11868, B0=>
      nx11876, B1=>nx11878);
   booth_integrtaion_4_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_31, QB=>nx11876, D=>nx5891, CLK=>clk, 
      R=>rst);
   ix11886 : inv01 port map ( Y=>nx11885, A=>weight_4(14));
   ix11889 : aoi22 port map ( Y=>nx11888, A0=>weight_4(15), A1=>nx5032, B0=>
      nx5036, B1=>nx5384);
   ix5385 : xnor2 port map ( Y=>nx5384, A0=>weight_4(15), A1=>nx5368);
   ix5369 : nor02ii port map ( Y=>nx5368, A0=>weight_4(14), A1=>nx5344);
   ix5379 : oai32 port map ( Y=>nx5378, A0=>nx11893, A1=>nx14512, A2=>nx5368, 
      B0=>nx11885, B1=>nx14516);
   ix11894 : nor02ii port map ( Y=>nx11893, A0=>nx5344, A1=>weight_4(14));
   ix5331 : oai32 port map ( Y=>nx5330, A0=>nx11897, A1=>nx14514, A2=>nx5320, 
      B0=>nx11849, B1=>nx14518);
   ix11898 : nor02ii port map ( Y=>nx11897, A0=>nx5296, A1=>weight_4(12));
   ix5283 : oai32 port map ( Y=>nx5282, A0=>nx11901, A1=>nx14514, A2=>nx5272, 
      B0=>nx11813, B1=>nx14518);
   ix11902 : nor02ii port map ( Y=>nx11901, A0=>nx5248, A1=>weight_4(10));
   ix5235 : oai32 port map ( Y=>nx5234, A0=>nx11905, A1=>nx14514, A2=>nx5224, 
      B0=>nx11777, B1=>nx14518);
   ix11906 : nor02ii port map ( Y=>nx11905, A0=>nx5200, A1=>weight_4(8));
   ix5187 : oai32 port map ( Y=>nx5186, A0=>nx11909, A1=>nx14514, A2=>nx5176, 
      B0=>nx11741, B1=>nx14518);
   ix11910 : nor02ii port map ( Y=>nx11909, A0=>nx5152, A1=>weight_4(6));
   ix5139 : oai32 port map ( Y=>nx5138, A0=>nx11913, A1=>nx14514, A2=>nx5128, 
      B0=>nx11705, B1=>nx14518);
   ix11914 : nor02ii port map ( Y=>nx11913, A0=>nx5104, A1=>weight_4(4));
   ix11917 : aoi32 port map ( Y=>nx11916, A0=>nx5050, A1=>nx5036, A2=>
      nx11649, B0=>weight_4(1), B1=>nx5032);
   booth_integrtaion_4_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_4_booth_output_16, QB=>nx11630, D=>nx6031, CLK=>clk, 
      R=>rst);
   booth_integrtaion_4_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_4_15, QB=>nx11920, D=>nx6041, CLK=>clk, R=>
      rst);
   ix5915 : xor2 port map ( Y=>label_4(1), A0=>nx11937, A1=>nx11939);
   ix11938 : nand02 port map ( Y=>nx11937, A0=>adderInput_4(0), A1=>
      booth_integration_output_4_0);
   ix11940 : xnor2 port map ( Y=>nx11939, A0=>booth_integration_output_4_1, 
      A1=>adderInput_4(1));
   ix5913 : xor2 port map ( Y=>label_4(2), A0=>nx11942, A1=>nx11945);
   ix11943 : aoi32 port map ( Y=>nx11942, A0=>adderInput_4(0), A1=>
      booth_integration_output_4_0, A2=>nx5772, B0=>adderInput_4(1), B1=>
      booth_integration_output_4_1);
   ix5911 : xnor2 port map ( Y=>label_4(3), A0=>nx5786, A1=>nx11951);
   ix5787 : oai22 port map ( Y=>nx5786, A0=>nx11942, A1=>nx11945, B0=>
      nx11949, B1=>nx11934);
   ix11950 : inv01 port map ( Y=>nx11949, A=>adderInput_4(2));
   ix11952 : xnor2 port map ( Y=>nx11951, A0=>booth_integration_output_4_3, 
      A1=>adderInput_4(3));
   ix5909 : xor2 port map ( Y=>label_4(4), A0=>nx11954, A1=>nx11957);
   ix11955 : aoi22 port map ( Y=>nx11954, A0=>adderInput_4(3), A1=>
      booth_integration_output_4_3, B0=>nx5786, B1=>nx5788);
   ix5907 : xnor2 port map ( Y=>label_4(5), A0=>nx5802, A1=>nx11963);
   ix5803 : oai22 port map ( Y=>nx5802, A0=>nx11954, A1=>nx11957, B0=>
      nx11961, B1=>nx11932);
   ix11962 : inv01 port map ( Y=>nx11961, A=>adderInput_4(4));
   ix11964 : xnor2 port map ( Y=>nx11963, A0=>booth_integration_output_4_5, 
      A1=>adderInput_4(5));
   ix5905 : xor2 port map ( Y=>label_4(6), A0=>nx11966, A1=>nx11969);
   ix11967 : aoi22 port map ( Y=>nx11966, A0=>adderInput_4(5), A1=>
      booth_integration_output_4_5, B0=>nx5802, B1=>nx5804);
   ix5903 : xnor2 port map ( Y=>label_4(7), A0=>nx5818, A1=>nx11975);
   ix5819 : oai22 port map ( Y=>nx5818, A0=>nx11966, A1=>nx11969, B0=>
      nx11973, B1=>nx11930);
   ix11974 : inv01 port map ( Y=>nx11973, A=>adderInput_4(6));
   ix11976 : xnor2 port map ( Y=>nx11975, A0=>booth_integration_output_4_7, 
      A1=>adderInput_4(7));
   ix5901 : xor2 port map ( Y=>label_4(8), A0=>nx11978, A1=>nx11981);
   ix11979 : aoi22 port map ( Y=>nx11978, A0=>adderInput_4(7), A1=>
      booth_integration_output_4_7, B0=>nx5818, B1=>nx5820);
   ix5899 : xnor2 port map ( Y=>label_4(9), A0=>nx5834, A1=>nx11987);
   ix5835 : oai22 port map ( Y=>nx5834, A0=>nx11978, A1=>nx11981, B0=>
      nx11985, B1=>nx11928);
   ix11986 : inv01 port map ( Y=>nx11985, A=>adderInput_4(8));
   ix11988 : xnor2 port map ( Y=>nx11987, A0=>booth_integration_output_4_9, 
      A1=>adderInput_4(9));
   ix5897 : xor2 port map ( Y=>label_4(10), A0=>nx11990, A1=>nx11993);
   ix11991 : aoi22 port map ( Y=>nx11990, A0=>adderInput_4(9), A1=>
      booth_integration_output_4_9, B0=>nx5834, B1=>nx5836);
   ix5895 : xnor2 port map ( Y=>label_4(11), A0=>nx5850, A1=>nx11999);
   ix5851 : oai22 port map ( Y=>nx5850, A0=>nx11990, A1=>nx11993, B0=>
      nx11997, B1=>nx11926);
   ix11998 : inv01 port map ( Y=>nx11997, A=>adderInput_4(10));
   ix12000 : xnor2 port map ( Y=>nx11999, A0=>booth_integration_output_4_11, 
      A1=>adderInput_4(11));
   ix5893 : xor2 port map ( Y=>label_4(12), A0=>nx12002, A1=>nx12005);
   ix12003 : aoi22 port map ( Y=>nx12002, A0=>adderInput_4(11), A1=>
      booth_integration_output_4_11, B0=>nx5850, B1=>nx5852);
   ix5891 : xnor2 port map ( Y=>label_4(13), A0=>nx5866, A1=>nx12011);
   ix5867 : oai22 port map ( Y=>nx5866, A0=>nx12002, A1=>nx12005, B0=>
      nx12009, B1=>nx11924);
   ix12010 : inv01 port map ( Y=>nx12009, A=>adderInput_4(12));
   ix12012 : xnor2 port map ( Y=>nx12011, A0=>booth_integration_output_4_13, 
      A1=>adderInput_4(13));
   ix5889 : xor2 port map ( Y=>label_4(14), A0=>nx12014, A1=>nx12017);
   ix12015 : aoi22 port map ( Y=>nx12014, A0=>adderInput_4(13), A1=>
      booth_integration_output_4_13, B0=>nx5866, B1=>nx5868);
   ix5887 : xnor2 port map ( Y=>label_4(15), A0=>nx5882, A1=>nx12023);
   ix5883 : oai22 port map ( Y=>nx5882, A0=>nx12014, A1=>nx12017, B0=>
      nx12021, B1=>nx11922);
   ix12022 : inv01 port map ( Y=>nx12021, A=>adderInput_4(14));
   booth_integrtaion_3_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_1, QB=>OPEN, D=>nx6711, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_2, QB=>nx12457, D=>nx6701, CLK=>clk, R=>rst
   );
   booth_integrtaion_3_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_3, QB=>OPEN, D=>nx6691, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_4, QB=>nx12455, D=>nx6681, CLK=>clk, R=>rst
   );
   booth_integrtaion_3_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_5, QB=>OPEN, D=>nx6671, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_6, QB=>nx12453, D=>nx6661, CLK=>clk, R=>rst
   );
   booth_integrtaion_3_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_7, QB=>OPEN, D=>nx6651, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_8, QB=>nx12451, D=>nx6641, CLK=>clk, R=>rst
   );
   booth_integrtaion_3_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_9, QB=>OPEN, D=>nx6631, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_10, QB=>nx12449, D=>nx6621, CLK=>clk, R=>
      rst);
   booth_integrtaion_3_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_11, QB=>OPEN, D=>nx6611, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_12, QB=>nx12447, D=>nx6601, CLK=>clk, R=>
      rst);
   booth_integrtaion_3_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_13, QB=>OPEN, D=>nx6591, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_14, QB=>nx12445, D=>nx6581, CLK=>clk, R=>
      rst);
   ix12075 : aoi22 port map ( Y=>nx12074, A0=>neuron(15), A1=>nx14306, B0=>
      nx6558, B1=>nx6564);
   booth_integrtaion_3_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_reg_output_0, QB=>OPEN, D=>nx6221, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_0, QB=>OPEN, D=>nx6207, CLK=>clk, 
      S=>nx14162);
   booth_integrtaion_3_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_reg_output_9, QB=>OPEN, D=>nx6401, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_9, QB=>OPEN, D=>nx6391, CLK=>clk, 
      R=>nx14162);
   booth_integrtaion_3_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_8, QB=>OPEN, D=>nx6381, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_8, QB=>OPEN, D=>nx6371, CLK=>clk, 
      R=>nx14162);
   booth_integrtaion_3_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_7, QB=>OPEN, D=>nx6361, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_7, QB=>OPEN, D=>nx6351, CLK=>clk, 
      R=>nx14162);
   booth_integrtaion_3_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_6, QB=>OPEN, D=>nx6341, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_6, QB=>OPEN, D=>nx6331, CLK=>clk, 
      R=>nx14162);
   booth_integrtaion_3_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_5, QB=>OPEN, D=>nx6321, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_5, QB=>OPEN, D=>nx6311, CLK=>clk, 
      R=>nx14162);
   booth_integrtaion_3_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_4, QB=>OPEN, D=>nx6301, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_4, QB=>OPEN, D=>nx6291, CLK=>clk, 
      R=>nx14160);
   booth_integrtaion_3_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_3, QB=>OPEN, D=>nx6281, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_3, QB=>OPEN, D=>nx6271, CLK=>clk, 
      R=>nx14160);
   booth_integrtaion_3_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_2, QB=>OPEN, D=>nx6261, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_2, QB=>OPEN, D=>nx6251, CLK=>clk, 
      R=>nx14160);
   booth_integrtaion_3_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_output_1, QB=>OPEN, D=>nx6241, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_3_shift_Reg_count_1, QB=>OPEN, D=>nx6231, CLK=>clk, 
      R=>nx14160);
   ix6202 : nand02 port map ( Y=>nx6201, A0=>nx14636, A1=>nx14292);
   booth_integrtaion_3_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx12121, D=>nx6201, CLK=>clk, S=>nx14160);
   ix6559 : nand02 port map ( Y=>nx6558, A0=>nx12142, A1=>nx12153);
   ix12143 : oai21 port map ( Y=>nx12142, A0=>nx6022, A1=>nx6018, B0=>
      weight_3(0));
   ix6412 : oai21 port map ( Y=>nx6411, A0=>nx12147, A1=>nx14520, B0=>
      nx12149);
   booth_integrtaion_3_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12147, D=>nx6411, CLK=>clk, R=>rst);
   booth_integrtaion_3_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_0, QB=>nx12026, D=>nx6721, CLK=>clk, R=>rst
   );
   ix12158 : xnor2 port map ( Y=>nx12157, A0=>nx6028, A1=>nx2954);
   ix6552 : oai21 port map ( Y=>nx6551, A0=>nx12163, A1=>nx14520, B0=>
      nx12165);
   booth_integrtaion_3_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_17, QB=>nx12163, D=>nx6551, CLK=>clk, 
      R=>rst);
   ix12166 : nand03 port map ( Y=>nx12165, A0=>nx14528, A1=>nx6536, A2=>
      nx14754);
   ix6537 : xnor2 port map ( Y=>nx6536, A0=>nx12168, A1=>nx2955);
   ix12169 : aoi22 port map ( Y=>nx12168, A0=>
      booth_integrtaion_3_booth_output_17, A1=>nx6052, B0=>nx6028, B1=>
      nx2954);
   ix6037 : nand02 port map ( Y=>nx6036, A0=>weight_3(1), A1=>weight_3(0));
   ix12173 : or02 port map ( Y=>nx12172, A0=>weight_3(0), A1=>weight_3(1));
   ix6542 : oai21 port map ( Y=>nx6541, A0=>nx12177, A1=>nx14520, B0=>
      nx12179);
   booth_integrtaion_3_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12177, D=>nx6541, CLK=>clk, R=>rst);
   ix12180 : nand03 port map ( Y=>nx12179, A0=>nx14528, A1=>nx6524, A2=>
      nx14754);
   ix6525 : xnor2 port map ( Y=>nx6524, A0=>nx6080, A1=>nx12190);
   ix6081 : oai22 port map ( Y=>nx6080, A0=>nx12168, A1=>nx12183, B0=>
      nx12177, B1=>nx14532);
   ix12186 : aoi32 port map ( Y=>nx12185, A0=>nx6062, A1=>nx6022, A2=>
      nx12188, B0=>weight_3(2), B1=>nx6018);
   ix6063 : oai21 port map ( Y=>nx6062, A0=>weight_3(0), A1=>weight_3(1), B0
      =>weight_3(2));
   ix12191 : xnor2 port map ( Y=>nx12190, A0=>
      booth_integrtaion_3_booth_output_19, A1=>nx6100);
   booth_integrtaion_3_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_19, QB=>OPEN, D=>nx6531, CLK=>clk, R
      =>rst);
   ix12196 : xnor2 port map ( Y=>nx12195, A0=>nx12197, A1=>nx12211);
   ix12198 : aoi22 port map ( Y=>nx12197, A0=>
      booth_integrtaion_3_booth_output_19, A1=>nx6100, B0=>nx6080, B1=>
      nx2956);
   ix6101 : oai32 port map ( Y=>nx6100, A0=>nx12200, A1=>nx14534, A2=>nx6090, 
      B0=>nx12206, B1=>nx14538);
   ix12201 : nor02ii port map ( Y=>nx12200, A0=>nx6066, A1=>weight_3(3));
   ix6067 : nor03_2x port map ( Y=>nx6066, A0=>weight_3(2), A1=>weight_3(0), 
      A2=>weight_3(1));
   ix6091 : nor04 port map ( Y=>nx6090, A0=>weight_3(3), A1=>weight_3(2), A2
      =>weight_3(0), A3=>weight_3(1));
   ix12207 : inv01 port map ( Y=>nx12206, A=>weight_3(3));
   ix6522 : oai21 port map ( Y=>nx6521, A0=>nx12215, A1=>nx14520, B0=>
      nx12217);
   booth_integrtaion_3_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12215, D=>nx6521, CLK=>clk, R=>rst);
   ix12218 : nand03 port map ( Y=>nx12217, A0=>nx14528, A1=>nx6500, A2=>
      nx14754);
   ix6501 : xnor2 port map ( Y=>nx6500, A0=>nx6128, A1=>nx12230);
   ix6129 : oai22 port map ( Y=>nx6128, A0=>nx12197, A1=>nx12211, B0=>
      nx12215, B1=>nx12221);
   ix12229 : inv01 port map ( Y=>nx12228, A=>weight_3(4));
   ix12231 : xnor2 port map ( Y=>nx12230, A0=>
      booth_integrtaion_3_booth_output_21, A1=>nx6148);
   booth_integrtaion_3_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_21, QB=>OPEN, D=>nx6511, CLK=>clk, R
      =>rst);
   ix12236 : xnor2 port map ( Y=>nx12235, A0=>nx12237, A1=>nx12247);
   ix12238 : aoi22 port map ( Y=>nx12237, A0=>
      booth_integrtaion_3_booth_output_21, A1=>nx6148, B0=>nx6128, B1=>
      nx2959);
   ix6149 : oai32 port map ( Y=>nx6148, A0=>nx12240, A1=>nx14534, A2=>nx6138, 
      B0=>nx12244, B1=>nx14538);
   ix12241 : nor02ii port map ( Y=>nx12240, A0=>nx6114, A1=>weight_3(5));
   ix6115 : nor02ii port map ( Y=>nx6114, A0=>weight_3(4), A1=>nx6090);
   ix6139 : nor02ii port map ( Y=>nx6138, A0=>weight_3(5), A1=>nx6114);
   ix12245 : inv01 port map ( Y=>nx12244, A=>weight_3(5));
   ix6502 : oai21 port map ( Y=>nx6501, A0=>nx12251, A1=>nx14520, B0=>
      nx12253);
   booth_integrtaion_3_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12251, D=>nx6501, CLK=>clk, R=>rst);
   ix12254 : nand03 port map ( Y=>nx12253, A0=>nx14528, A1=>nx6476, A2=>
      nx14522);
   ix6477 : xnor2 port map ( Y=>nx6476, A0=>nx6176, A1=>nx12266);
   ix6177 : oai22 port map ( Y=>nx6176, A0=>nx12237, A1=>nx12247, B0=>
      nx12251, B1=>nx12257);
   ix12265 : inv01 port map ( Y=>nx12264, A=>weight_3(6));
   ix12267 : xnor2 port map ( Y=>nx12266, A0=>
      booth_integrtaion_3_booth_output_23, A1=>nx6196);
   booth_integrtaion_3_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_23, QB=>OPEN, D=>nx6491, CLK=>clk, R
      =>rst);
   ix12272 : xnor2 port map ( Y=>nx12271, A0=>nx12273, A1=>nx12283);
   ix12274 : aoi22 port map ( Y=>nx12273, A0=>
      booth_integrtaion_3_booth_output_23, A1=>nx6196, B0=>nx6176, B1=>
      nx2961);
   ix6197 : oai32 port map ( Y=>nx6196, A0=>nx12276, A1=>nx14534, A2=>nx6186, 
      B0=>nx12280, B1=>nx14538);
   ix12277 : nor02ii port map ( Y=>nx12276, A0=>nx6162, A1=>weight_3(7));
   ix6163 : nor02ii port map ( Y=>nx6162, A0=>weight_3(6), A1=>nx6138);
   ix6187 : nor02ii port map ( Y=>nx6186, A0=>weight_3(7), A1=>nx6162);
   ix12281 : inv01 port map ( Y=>nx12280, A=>weight_3(7));
   ix6482 : oai21 port map ( Y=>nx6481, A0=>nx12287, A1=>nx14522, B0=>
      nx12289);
   booth_integrtaion_3_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12287, D=>nx6481, CLK=>clk, R=>rst);
   ix12290 : nand03 port map ( Y=>nx12289, A0=>nx14528, A1=>nx6452, A2=>
      nx14522);
   ix6453 : xnor2 port map ( Y=>nx6452, A0=>nx6224, A1=>nx12302);
   ix6225 : oai22 port map ( Y=>nx6224, A0=>nx12273, A1=>nx12283, B0=>
      nx12287, B1=>nx12293);
   ix12301 : inv01 port map ( Y=>nx12300, A=>weight_3(8));
   ix12303 : xnor2 port map ( Y=>nx12302, A0=>
      booth_integrtaion_3_booth_output_25, A1=>nx6244);
   booth_integrtaion_3_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_25, QB=>OPEN, D=>nx6471, CLK=>clk, R
      =>rst);
   ix12308 : xnor2 port map ( Y=>nx12307, A0=>nx12309, A1=>nx12319);
   ix12310 : aoi22 port map ( Y=>nx12309, A0=>
      booth_integrtaion_3_booth_output_25, A1=>nx6244, B0=>nx6224, B1=>
      nx2963);
   ix6245 : oai32 port map ( Y=>nx6244, A0=>nx12312, A1=>nx14534, A2=>nx6234, 
      B0=>nx12316, B1=>nx14538);
   ix12313 : nor02ii port map ( Y=>nx12312, A0=>nx6210, A1=>weight_3(9));
   ix6211 : nor02ii port map ( Y=>nx6210, A0=>weight_3(8), A1=>nx6186);
   ix6235 : nor02ii port map ( Y=>nx6234, A0=>weight_3(9), A1=>nx6210);
   ix12317 : inv01 port map ( Y=>nx12316, A=>weight_3(9));
   ix6462 : oai21 port map ( Y=>nx6461, A0=>nx12323, A1=>nx14522, B0=>
      nx12325);
   booth_integrtaion_3_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12323, D=>nx6461, CLK=>clk, R=>rst);
   ix12326 : nand03 port map ( Y=>nx12325, A0=>nx14528, A1=>nx6428, A2=>
      nx14522);
   ix6429 : xnor2 port map ( Y=>nx6428, A0=>nx6272, A1=>nx12338);
   ix6273 : oai22 port map ( Y=>nx6272, A0=>nx12309, A1=>nx12319, B0=>
      nx12323, B1=>nx12329);
   ix12337 : inv01 port map ( Y=>nx12336, A=>weight_3(10));
   ix12339 : xnor2 port map ( Y=>nx12338, A0=>
      booth_integrtaion_3_booth_output_27, A1=>nx6292);
   booth_integrtaion_3_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_27, QB=>OPEN, D=>nx6451, CLK=>clk, R
      =>rst);
   ix12344 : xnor2 port map ( Y=>nx12343, A0=>nx12345, A1=>nx12355);
   ix12346 : aoi22 port map ( Y=>nx12345, A0=>
      booth_integrtaion_3_booth_output_27, A1=>nx6292, B0=>nx6272, B1=>
      nx2965);
   ix6293 : oai32 port map ( Y=>nx6292, A0=>nx12348, A1=>nx14534, A2=>nx6282, 
      B0=>nx12352, B1=>nx14538);
   ix12349 : nor02ii port map ( Y=>nx12348, A0=>nx6258, A1=>weight_3(11));
   ix6259 : nor02ii port map ( Y=>nx6258, A0=>weight_3(10), A1=>nx6234);
   ix6283 : nor02ii port map ( Y=>nx6282, A0=>weight_3(11), A1=>nx6258);
   ix12353 : inv01 port map ( Y=>nx12352, A=>weight_3(11));
   ix6442 : oai21 port map ( Y=>nx6441, A0=>nx12359, A1=>nx14522, B0=>
      nx12361);
   booth_integrtaion_3_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12359, D=>nx6441, CLK=>clk, R=>rst);
   ix12362 : nand03 port map ( Y=>nx12361, A0=>nx14762, A1=>nx6404, A2=>
      nx14522);
   ix6405 : xnor2 port map ( Y=>nx6404, A0=>nx6320, A1=>nx12374);
   ix6321 : oai22 port map ( Y=>nx6320, A0=>nx12345, A1=>nx12355, B0=>
      nx12359, B1=>nx12365);
   ix12373 : inv01 port map ( Y=>nx12372, A=>weight_3(12));
   ix12375 : xnor2 port map ( Y=>nx12374, A0=>
      booth_integrtaion_3_booth_output_29, A1=>nx6340);
   booth_integrtaion_3_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_29, QB=>OPEN, D=>nx6431, CLK=>clk, R
      =>rst);
   ix12380 : xnor2 port map ( Y=>nx12379, A0=>nx12381, A1=>nx12391);
   ix12382 : aoi22 port map ( Y=>nx12381, A0=>
      booth_integrtaion_3_booth_output_29, A1=>nx6340, B0=>nx6320, B1=>
      nx2967);
   ix6341 : oai32 port map ( Y=>nx6340, A0=>nx12384, A1=>nx14534, A2=>nx6330, 
      B0=>nx12388, B1=>nx14538);
   ix12385 : nor02ii port map ( Y=>nx12384, A0=>nx6306, A1=>weight_3(13));
   ix6307 : nor02ii port map ( Y=>nx6306, A0=>weight_3(12), A1=>nx6282);
   ix6331 : nor02ii port map ( Y=>nx6330, A0=>weight_3(13), A1=>nx6306);
   ix12389 : inv01 port map ( Y=>nx12388, A=>weight_3(13));
   ix12397 : xnor2 port map ( Y=>nx12396, A0=>nx6368, A1=>nx6378);
   ix6369 : oai22 port map ( Y=>nx6368, A0=>nx12381, A1=>nx12391, B0=>
      nx12399, B1=>nx12401);
   booth_integrtaion_3_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_31, QB=>nx12399, D=>nx6421, CLK=>clk, 
      R=>rst);
   ix12409 : inv01 port map ( Y=>nx12408, A=>weight_3(14));
   ix12412 : aoi22 port map ( Y=>nx12411, A0=>weight_3(15), A1=>nx6018, B0=>
      nx6022, B1=>nx6370);
   ix6371 : xnor2 port map ( Y=>nx6370, A0=>weight_3(15), A1=>nx6354);
   ix6355 : nor02ii port map ( Y=>nx6354, A0=>weight_3(14), A1=>nx6330);
   ix6365 : oai32 port map ( Y=>nx6364, A0=>nx12416, A1=>nx14534, A2=>nx6354, 
      B0=>nx12408, B1=>nx14538);
   ix12417 : nor02ii port map ( Y=>nx12416, A0=>nx6330, A1=>weight_3(14));
   ix6317 : oai32 port map ( Y=>nx6316, A0=>nx12420, A1=>nx14536, A2=>nx6306, 
      B0=>nx12372, B1=>nx14540);
   ix12421 : nor02ii port map ( Y=>nx12420, A0=>nx6282, A1=>weight_3(12));
   ix6269 : oai32 port map ( Y=>nx6268, A0=>nx12424, A1=>nx14536, A2=>nx6258, 
      B0=>nx12336, B1=>nx14540);
   ix12425 : nor02ii port map ( Y=>nx12424, A0=>nx6234, A1=>weight_3(10));
   ix6221 : oai32 port map ( Y=>nx6220, A0=>nx12428, A1=>nx14536, A2=>nx6210, 
      B0=>nx12300, B1=>nx14540);
   ix12429 : nor02ii port map ( Y=>nx12428, A0=>nx6186, A1=>weight_3(8));
   ix6173 : oai32 port map ( Y=>nx6172, A0=>nx12432, A1=>nx14536, A2=>nx6162, 
      B0=>nx12264, B1=>nx14540);
   ix12433 : nor02ii port map ( Y=>nx12432, A0=>nx6138, A1=>weight_3(6));
   ix6125 : oai32 port map ( Y=>nx6124, A0=>nx12436, A1=>nx14536, A2=>nx6114, 
      B0=>nx12228, B1=>nx14540);
   ix12437 : nor02ii port map ( Y=>nx12436, A0=>nx6090, A1=>weight_3(4));
   ix12440 : aoi32 port map ( Y=>nx12439, A0=>nx6036, A1=>nx6022, A2=>
      nx12172, B0=>weight_3(1), B1=>nx6018);
   booth_integrtaion_3_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_3_booth_output_16, QB=>nx12153, D=>nx6561, CLK=>clk, 
      R=>rst);
   booth_integrtaion_3_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_3_15, QB=>nx12443, D=>nx6571, CLK=>clk, R=>
      rst);
   ix6901 : xor2 port map ( Y=>label_3(1), A0=>nx12460, A1=>nx12462);
   ix12461 : nand02 port map ( Y=>nx12460, A0=>adderInput_3(0), A1=>
      booth_integration_output_3_0);
   ix12463 : xnor2 port map ( Y=>nx12462, A0=>booth_integration_output_3_1, 
      A1=>adderInput_3(1));
   ix6899 : xor2 port map ( Y=>label_3(2), A0=>nx12465, A1=>nx12468);
   ix12466 : aoi32 port map ( Y=>nx12465, A0=>adderInput_3(0), A1=>
      booth_integration_output_3_0, A2=>nx6758, B0=>adderInput_3(1), B1=>
      booth_integration_output_3_1);
   ix6897 : xnor2 port map ( Y=>label_3(3), A0=>nx6772, A1=>nx12474);
   ix6773 : oai22 port map ( Y=>nx6772, A0=>nx12465, A1=>nx12468, B0=>
      nx12472, B1=>nx12457);
   ix12473 : inv01 port map ( Y=>nx12472, A=>adderInput_3(2));
   ix12475 : xnor2 port map ( Y=>nx12474, A0=>booth_integration_output_3_3, 
      A1=>adderInput_3(3));
   ix6895 : xor2 port map ( Y=>label_3(4), A0=>nx12477, A1=>nx12480);
   ix12478 : aoi22 port map ( Y=>nx12477, A0=>adderInput_3(3), A1=>
      booth_integration_output_3_3, B0=>nx6772, B1=>nx6774);
   ix6893 : xnor2 port map ( Y=>label_3(5), A0=>nx6788, A1=>nx12486);
   ix6789 : oai22 port map ( Y=>nx6788, A0=>nx12477, A1=>nx12480, B0=>
      nx12484, B1=>nx12455);
   ix12485 : inv01 port map ( Y=>nx12484, A=>adderInput_3(4));
   ix12487 : xnor2 port map ( Y=>nx12486, A0=>booth_integration_output_3_5, 
      A1=>adderInput_3(5));
   ix6891 : xor2 port map ( Y=>label_3(6), A0=>nx12489, A1=>nx12492);
   ix12490 : aoi22 port map ( Y=>nx12489, A0=>adderInput_3(5), A1=>
      booth_integration_output_3_5, B0=>nx6788, B1=>nx6790);
   ix6889 : xnor2 port map ( Y=>label_3(7), A0=>nx6804, A1=>nx12498);
   ix6805 : oai22 port map ( Y=>nx6804, A0=>nx12489, A1=>nx12492, B0=>
      nx12496, B1=>nx12453);
   ix12497 : inv01 port map ( Y=>nx12496, A=>adderInput_3(6));
   ix12499 : xnor2 port map ( Y=>nx12498, A0=>booth_integration_output_3_7, 
      A1=>adderInput_3(7));
   ix6887 : xor2 port map ( Y=>label_3(8), A0=>nx12501, A1=>nx12504);
   ix12502 : aoi22 port map ( Y=>nx12501, A0=>adderInput_3(7), A1=>
      booth_integration_output_3_7, B0=>nx6804, B1=>nx6806);
   ix6885 : xnor2 port map ( Y=>label_3(9), A0=>nx6820, A1=>nx12510);
   ix6821 : oai22 port map ( Y=>nx6820, A0=>nx12501, A1=>nx12504, B0=>
      nx12508, B1=>nx12451);
   ix12509 : inv01 port map ( Y=>nx12508, A=>adderInput_3(8));
   ix12511 : xnor2 port map ( Y=>nx12510, A0=>booth_integration_output_3_9, 
      A1=>adderInput_3(9));
   ix6883 : xor2 port map ( Y=>label_3(10), A0=>nx12513, A1=>nx12516);
   ix12514 : aoi22 port map ( Y=>nx12513, A0=>adderInput_3(9), A1=>
      booth_integration_output_3_9, B0=>nx6820, B1=>nx6822);
   ix6881 : xnor2 port map ( Y=>label_3(11), A0=>nx6836, A1=>nx12522);
   ix6837 : oai22 port map ( Y=>nx6836, A0=>nx12513, A1=>nx12516, B0=>
      nx12520, B1=>nx12449);
   ix12521 : inv01 port map ( Y=>nx12520, A=>adderInput_3(10));
   ix12523 : xnor2 port map ( Y=>nx12522, A0=>booth_integration_output_3_11, 
      A1=>adderInput_3(11));
   ix6879 : xor2 port map ( Y=>label_3(12), A0=>nx12525, A1=>nx12528);
   ix12526 : aoi22 port map ( Y=>nx12525, A0=>adderInput_3(11), A1=>
      booth_integration_output_3_11, B0=>nx6836, B1=>nx6838);
   ix6877 : xnor2 port map ( Y=>label_3(13), A0=>nx6852, A1=>nx12534);
   ix6853 : oai22 port map ( Y=>nx6852, A0=>nx12525, A1=>nx12528, B0=>
      nx12532, B1=>nx12447);
   ix12533 : inv01 port map ( Y=>nx12532, A=>adderInput_3(12));
   ix12535 : xnor2 port map ( Y=>nx12534, A0=>booth_integration_output_3_13, 
      A1=>adderInput_3(13));
   ix6875 : xor2 port map ( Y=>label_3(14), A0=>nx12537, A1=>nx12540);
   ix12538 : aoi22 port map ( Y=>nx12537, A0=>adderInput_3(13), A1=>
      booth_integration_output_3_13, B0=>nx6852, B1=>nx6854);
   ix6873 : xnor2 port map ( Y=>label_3(15), A0=>nx6868, A1=>nx12546);
   ix6869 : oai22 port map ( Y=>nx6868, A0=>nx12537, A1=>nx12540, B0=>
      nx12544, B1=>nx12445);
   ix12545 : inv01 port map ( Y=>nx12544, A=>adderInput_3(14));
   booth_integrtaion_2_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_1, QB=>OPEN, D=>nx7241, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_2, QB=>nx12980, D=>nx7231, CLK=>clk, R=>rst
   );
   booth_integrtaion_2_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_3, QB=>OPEN, D=>nx7221, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_4, QB=>nx12978, D=>nx7211, CLK=>clk, R=>rst
   );
   booth_integrtaion_2_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_5, QB=>OPEN, D=>nx7201, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_6, QB=>nx12976, D=>nx7191, CLK=>clk, R=>rst
   );
   booth_integrtaion_2_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_7, QB=>OPEN, D=>nx7181, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_8, QB=>nx12974, D=>nx7171, CLK=>clk, R=>rst
   );
   booth_integrtaion_2_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_9, QB=>OPEN, D=>nx7161, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_10, QB=>nx12972, D=>nx7151, CLK=>clk, R=>
      rst);
   booth_integrtaion_2_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_11, QB=>OPEN, D=>nx7141, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_12, QB=>nx12970, D=>nx7131, CLK=>clk, R=>
      rst);
   booth_integrtaion_2_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_13, QB=>OPEN, D=>nx7121, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_14, QB=>nx12968, D=>nx7111, CLK=>clk, R=>
      rst);
   ix12598 : aoi22 port map ( Y=>nx12597, A0=>neuron(15), A1=>nx14328, B0=>
      nx7544, B1=>nx7550);
   booth_integrtaion_2_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_reg_output_0, QB=>OPEN, D=>nx6751, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_0, QB=>OPEN, D=>nx6737, CLK=>clk, 
      S=>nx14166);
   booth_integrtaion_2_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_reg_output_9, QB=>OPEN, D=>nx6931, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_9, QB=>OPEN, D=>nx6921, CLK=>clk, 
      R=>nx14166);
   booth_integrtaion_2_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_8, QB=>OPEN, D=>nx6911, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_8, QB=>OPEN, D=>nx6901, CLK=>clk, 
      R=>nx14166);
   booth_integrtaion_2_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_7, QB=>OPEN, D=>nx6891, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_7, QB=>OPEN, D=>nx6881, CLK=>clk, 
      R=>nx14164);
   booth_integrtaion_2_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_6, QB=>OPEN, D=>nx6871, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_6, QB=>OPEN, D=>nx6861, CLK=>clk, 
      R=>nx14164);
   booth_integrtaion_2_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_5, QB=>OPEN, D=>nx6851, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_5, QB=>OPEN, D=>nx6841, CLK=>clk, 
      R=>nx14164);
   booth_integrtaion_2_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_4, QB=>OPEN, D=>nx6831, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_4, QB=>OPEN, D=>nx6821, CLK=>clk, 
      R=>nx14164);
   booth_integrtaion_2_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_3, QB=>OPEN, D=>nx6811, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_3, QB=>OPEN, D=>nx6801, CLK=>clk, 
      R=>nx14164);
   booth_integrtaion_2_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_2, QB=>OPEN, D=>nx6791, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_2, QB=>OPEN, D=>nx6781, CLK=>clk, 
      R=>nx14164);
   booth_integrtaion_2_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_output_1, QB=>OPEN, D=>nx6771, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_2_shift_Reg_count_1, QB=>OPEN, D=>nx6761, CLK=>clk, 
      R=>nx14162);
   ix6732 : nand02 port map ( Y=>nx6731, A0=>nx14640, A1=>nx14314);
   booth_integrtaion_2_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx12644, D=>nx6731, CLK=>clk, S=>nx14164);
   ix7545 : nand02 port map ( Y=>nx7544, A0=>nx12665, A1=>nx12676);
   ix12666 : oai21 port map ( Y=>nx12665, A0=>nx7008, A1=>nx7004, B0=>
      weight_2(0));
   ix6942 : oai21 port map ( Y=>nx6941, A0=>nx12670, A1=>nx14542, B0=>
      nx12672);
   booth_integrtaion_2_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12670, D=>nx6941, CLK=>clk, R=>rst);
   booth_integrtaion_2_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_0, QB=>nx12549, D=>nx7251, CLK=>clk, R=>rst
   );
   ix12681 : xnor2 port map ( Y=>nx12680, A0=>nx7014, A1=>nx2970);
   ix7082 : oai21 port map ( Y=>nx7081, A0=>nx12686, A1=>nx14542, B0=>
      nx12688);
   booth_integrtaion_2_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_17, QB=>nx12686, D=>nx7081, CLK=>clk, 
      R=>rst);
   ix12689 : nand03 port map ( Y=>nx12688, A0=>nx14550, A1=>nx7522, A2=>
      nx14770);
   ix7523 : xnor2 port map ( Y=>nx7522, A0=>nx12691, A1=>nx2971);
   ix12692 : aoi22 port map ( Y=>nx12691, A0=>
      booth_integrtaion_2_booth_output_17, A1=>nx7038, B0=>nx7014, B1=>
      nx2970);
   ix7023 : nand02 port map ( Y=>nx7022, A0=>weight_2(1), A1=>weight_2(0));
   ix12696 : or02 port map ( Y=>nx12695, A0=>weight_2(0), A1=>weight_2(1));
   ix7072 : oai21 port map ( Y=>nx7071, A0=>nx12700, A1=>nx14542, B0=>
      nx12702);
   booth_integrtaion_2_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12700, D=>nx7071, CLK=>clk, R=>rst);
   ix12703 : nand03 port map ( Y=>nx12702, A0=>nx14550, A1=>nx7510, A2=>
      nx14770);
   ix7511 : xnor2 port map ( Y=>nx7510, A0=>nx7066, A1=>nx12713);
   ix7067 : oai22 port map ( Y=>nx7066, A0=>nx12691, A1=>nx12706, B0=>
      nx12700, B1=>nx14554);
   ix12709 : aoi32 port map ( Y=>nx12708, A0=>nx7048, A1=>nx7008, A2=>
      nx12711, B0=>weight_2(2), B1=>nx7004);
   ix7049 : oai21 port map ( Y=>nx7048, A0=>weight_2(0), A1=>weight_2(1), B0
      =>weight_2(2));
   ix12714 : xnor2 port map ( Y=>nx12713, A0=>
      booth_integrtaion_2_booth_output_19, A1=>nx7086);
   booth_integrtaion_2_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_19, QB=>OPEN, D=>nx7061, CLK=>clk, R
      =>rst);
   ix12719 : xnor2 port map ( Y=>nx12718, A0=>nx12720, A1=>nx12734);
   ix12721 : aoi22 port map ( Y=>nx12720, A0=>
      booth_integrtaion_2_booth_output_19, A1=>nx7086, B0=>nx7066, B1=>
      nx2972);
   ix7087 : oai32 port map ( Y=>nx7086, A0=>nx12723, A1=>nx14556, A2=>nx7076, 
      B0=>nx12729, B1=>nx14560);
   ix12724 : nor02ii port map ( Y=>nx12723, A0=>nx7052, A1=>weight_2(3));
   ix7053 : nor03_2x port map ( Y=>nx7052, A0=>weight_2(2), A1=>weight_2(0), 
      A2=>weight_2(1));
   ix7077 : nor04 port map ( Y=>nx7076, A0=>weight_2(3), A1=>weight_2(2), A2
      =>weight_2(0), A3=>weight_2(1));
   ix12730 : inv01 port map ( Y=>nx12729, A=>weight_2(3));
   ix7052 : oai21 port map ( Y=>nx7051, A0=>nx12738, A1=>nx14542, B0=>
      nx12740);
   booth_integrtaion_2_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12738, D=>nx7051, CLK=>clk, R=>rst);
   ix12741 : nand03 port map ( Y=>nx12740, A0=>nx14550, A1=>nx7486, A2=>
      nx14770);
   ix7487 : xnor2 port map ( Y=>nx7486, A0=>nx7114, A1=>nx12753);
   ix7115 : oai22 port map ( Y=>nx7114, A0=>nx12720, A1=>nx12734, B0=>
      nx12738, B1=>nx12744);
   ix12752 : inv01 port map ( Y=>nx12751, A=>weight_2(4));
   ix12754 : xnor2 port map ( Y=>nx12753, A0=>
      booth_integrtaion_2_booth_output_21, A1=>nx7134);
   booth_integrtaion_2_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_21, QB=>OPEN, D=>nx7041, CLK=>clk, R
      =>rst);
   ix12759 : xnor2 port map ( Y=>nx12758, A0=>nx12760, A1=>nx12770);
   ix12761 : aoi22 port map ( Y=>nx12760, A0=>
      booth_integrtaion_2_booth_output_21, A1=>nx7134, B0=>nx7114, B1=>
      nx2974);
   ix7135 : oai32 port map ( Y=>nx7134, A0=>nx12763, A1=>nx14556, A2=>nx7124, 
      B0=>nx12767, B1=>nx14560);
   ix12764 : nor02ii port map ( Y=>nx12763, A0=>nx7100, A1=>weight_2(5));
   ix7101 : nor02ii port map ( Y=>nx7100, A0=>weight_2(4), A1=>nx7076);
   ix7125 : nor02ii port map ( Y=>nx7124, A0=>weight_2(5), A1=>nx7100);
   ix12768 : inv01 port map ( Y=>nx12767, A=>weight_2(5));
   ix7032 : oai21 port map ( Y=>nx7031, A0=>nx12774, A1=>nx14542, B0=>
      nx12776);
   booth_integrtaion_2_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12774, D=>nx7031, CLK=>clk, R=>rst);
   ix12777 : nand03 port map ( Y=>nx12776, A0=>nx14550, A1=>nx7462, A2=>
      nx14544);
   ix7463 : xnor2 port map ( Y=>nx7462, A0=>nx7162, A1=>nx12789);
   ix7163 : oai22 port map ( Y=>nx7162, A0=>nx12760, A1=>nx12770, B0=>
      nx12774, B1=>nx12780);
   ix12788 : inv01 port map ( Y=>nx12787, A=>weight_2(6));
   ix12790 : xnor2 port map ( Y=>nx12789, A0=>
      booth_integrtaion_2_booth_output_23, A1=>nx7182);
   booth_integrtaion_2_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_23, QB=>OPEN, D=>nx7021, CLK=>clk, R
      =>rst);
   ix12795 : xnor2 port map ( Y=>nx12794, A0=>nx12796, A1=>nx12806);
   ix12797 : aoi22 port map ( Y=>nx12796, A0=>
      booth_integrtaion_2_booth_output_23, A1=>nx7182, B0=>nx7162, B1=>
      nx2976);
   ix7183 : oai32 port map ( Y=>nx7182, A0=>nx12799, A1=>nx14556, A2=>nx7172, 
      B0=>nx12803, B1=>nx14560);
   ix12800 : nor02ii port map ( Y=>nx12799, A0=>nx7148, A1=>weight_2(7));
   ix7149 : nor02ii port map ( Y=>nx7148, A0=>weight_2(6), A1=>nx7124);
   ix7173 : nor02ii port map ( Y=>nx7172, A0=>weight_2(7), A1=>nx7148);
   ix12804 : inv01 port map ( Y=>nx12803, A=>weight_2(7));
   ix7012 : oai21 port map ( Y=>nx7011, A0=>nx12810, A1=>nx14544, B0=>
      nx12812);
   booth_integrtaion_2_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12810, D=>nx7011, CLK=>clk, R=>rst);
   ix12813 : nand03 port map ( Y=>nx12812, A0=>nx14550, A1=>nx7438, A2=>
      nx14544);
   ix7439 : xnor2 port map ( Y=>nx7438, A0=>nx7210, A1=>nx12825);
   ix7211 : oai22 port map ( Y=>nx7210, A0=>nx12796, A1=>nx12806, B0=>
      nx12810, B1=>nx12816);
   ix12824 : inv01 port map ( Y=>nx12823, A=>weight_2(8));
   ix12826 : xnor2 port map ( Y=>nx12825, A0=>
      booth_integrtaion_2_booth_output_25, A1=>nx7230);
   booth_integrtaion_2_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_25, QB=>OPEN, D=>nx7001, CLK=>clk, R
      =>rst);
   ix12831 : xnor2 port map ( Y=>nx12830, A0=>nx12832, A1=>nx12842);
   ix12833 : aoi22 port map ( Y=>nx12832, A0=>
      booth_integrtaion_2_booth_output_25, A1=>nx7230, B0=>nx7210, B1=>
      nx2978);
   ix7231 : oai32 port map ( Y=>nx7230, A0=>nx12835, A1=>nx14556, A2=>nx7220, 
      B0=>nx12839, B1=>nx14560);
   ix12836 : nor02ii port map ( Y=>nx12835, A0=>nx7196, A1=>weight_2(9));
   ix7197 : nor02ii port map ( Y=>nx7196, A0=>weight_2(8), A1=>nx7172);
   ix7221 : nor02ii port map ( Y=>nx7220, A0=>weight_2(9), A1=>nx7196);
   ix12840 : inv01 port map ( Y=>nx12839, A=>weight_2(9));
   ix6992 : oai21 port map ( Y=>nx6991, A0=>nx12846, A1=>nx14544, B0=>
      nx12848);
   booth_integrtaion_2_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12846, D=>nx6991, CLK=>clk, R=>rst);
   ix12849 : nand03 port map ( Y=>nx12848, A0=>nx14550, A1=>nx7414, A2=>
      nx14544);
   ix7415 : xnor2 port map ( Y=>nx7414, A0=>nx7258, A1=>nx12861);
   ix7259 : oai22 port map ( Y=>nx7258, A0=>nx12832, A1=>nx12842, B0=>
      nx12846, B1=>nx12852);
   ix12860 : inv01 port map ( Y=>nx12859, A=>weight_2(10));
   ix12862 : xnor2 port map ( Y=>nx12861, A0=>
      booth_integrtaion_2_booth_output_27, A1=>nx7278);
   booth_integrtaion_2_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_27, QB=>OPEN, D=>nx6981, CLK=>clk, R
      =>rst);
   ix12867 : xnor2 port map ( Y=>nx12866, A0=>nx12868, A1=>nx12878);
   ix12869 : aoi22 port map ( Y=>nx12868, A0=>
      booth_integrtaion_2_booth_output_27, A1=>nx7278, B0=>nx7258, B1=>
      nx2980);
   ix7279 : oai32 port map ( Y=>nx7278, A0=>nx12871, A1=>nx14556, A2=>nx7268, 
      B0=>nx12875, B1=>nx14560);
   ix12872 : nor02ii port map ( Y=>nx12871, A0=>nx7244, A1=>weight_2(11));
   ix7245 : nor02ii port map ( Y=>nx7244, A0=>weight_2(10), A1=>nx7220);
   ix7269 : nor02ii port map ( Y=>nx7268, A0=>weight_2(11), A1=>nx7244);
   ix12876 : inv01 port map ( Y=>nx12875, A=>weight_2(11));
   ix6972 : oai21 port map ( Y=>nx6971, A0=>nx12882, A1=>nx14544, B0=>
      nx12884);
   booth_integrtaion_2_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx12882, D=>nx6971, CLK=>clk, R=>rst);
   ix12885 : nand03 port map ( Y=>nx12884, A0=>nx14778, A1=>nx7390, A2=>
      nx14544);
   ix7391 : xnor2 port map ( Y=>nx7390, A0=>nx7306, A1=>nx12897);
   ix7307 : oai22 port map ( Y=>nx7306, A0=>nx12868, A1=>nx12878, B0=>
      nx12882, B1=>nx12888);
   ix12896 : inv01 port map ( Y=>nx12895, A=>weight_2(12));
   ix12898 : xnor2 port map ( Y=>nx12897, A0=>
      booth_integrtaion_2_booth_output_29, A1=>nx7326);
   booth_integrtaion_2_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_29, QB=>OPEN, D=>nx6961, CLK=>clk, R
      =>rst);
   ix12903 : xnor2 port map ( Y=>nx12902, A0=>nx12904, A1=>nx12914);
   ix12905 : aoi22 port map ( Y=>nx12904, A0=>
      booth_integrtaion_2_booth_output_29, A1=>nx7326, B0=>nx7306, B1=>
      nx2982);
   ix7327 : oai32 port map ( Y=>nx7326, A0=>nx12907, A1=>nx14556, A2=>nx7316, 
      B0=>nx12911, B1=>nx14560);
   ix12908 : nor02ii port map ( Y=>nx12907, A0=>nx7292, A1=>weight_2(13));
   ix7293 : nor02ii port map ( Y=>nx7292, A0=>weight_2(12), A1=>nx7268);
   ix7317 : nor02ii port map ( Y=>nx7316, A0=>weight_2(13), A1=>nx7292);
   ix12912 : inv01 port map ( Y=>nx12911, A=>weight_2(13));
   ix12920 : xnor2 port map ( Y=>nx12919, A0=>nx7354, A1=>nx7364);
   ix7355 : oai22 port map ( Y=>nx7354, A0=>nx12904, A1=>nx12914, B0=>
      nx12922, B1=>nx12924);
   booth_integrtaion_2_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_31, QB=>nx12922, D=>nx6951, CLK=>clk, 
      R=>rst);
   ix12932 : inv01 port map ( Y=>nx12931, A=>weight_2(14));
   ix12935 : aoi22 port map ( Y=>nx12934, A0=>weight_2(15), A1=>nx7004, B0=>
      nx7008, B1=>nx7356);
   ix7357 : xnor2 port map ( Y=>nx7356, A0=>weight_2(15), A1=>nx7340);
   ix7341 : nor02ii port map ( Y=>nx7340, A0=>weight_2(14), A1=>nx7316);
   ix7351 : oai32 port map ( Y=>nx7350, A0=>nx12939, A1=>nx14556, A2=>nx7340, 
      B0=>nx12931, B1=>nx14560);
   ix12940 : nor02ii port map ( Y=>nx12939, A0=>nx7316, A1=>weight_2(14));
   ix7303 : oai32 port map ( Y=>nx7302, A0=>nx12943, A1=>nx14558, A2=>nx7292, 
      B0=>nx12895, B1=>nx14562);
   ix12944 : nor02ii port map ( Y=>nx12943, A0=>nx7268, A1=>weight_2(12));
   ix7255 : oai32 port map ( Y=>nx7254, A0=>nx12947, A1=>nx14558, A2=>nx7244, 
      B0=>nx12859, B1=>nx14562);
   ix12948 : nor02ii port map ( Y=>nx12947, A0=>nx7220, A1=>weight_2(10));
   ix7207 : oai32 port map ( Y=>nx7206, A0=>nx12951, A1=>nx14558, A2=>nx7196, 
      B0=>nx12823, B1=>nx14562);
   ix12952 : nor02ii port map ( Y=>nx12951, A0=>nx7172, A1=>weight_2(8));
   ix7159 : oai32 port map ( Y=>nx7158, A0=>nx12955, A1=>nx14558, A2=>nx7148, 
      B0=>nx12787, B1=>nx14562);
   ix12956 : nor02ii port map ( Y=>nx12955, A0=>nx7124, A1=>weight_2(6));
   ix7111 : oai32 port map ( Y=>nx7110, A0=>nx12959, A1=>nx14558, A2=>nx7100, 
      B0=>nx12751, B1=>nx14562);
   ix12960 : nor02ii port map ( Y=>nx12959, A0=>nx7076, A1=>weight_2(4));
   ix12963 : aoi32 port map ( Y=>nx12962, A0=>nx7022, A1=>nx7008, A2=>
      nx12695, B0=>weight_2(1), B1=>nx7004);
   booth_integrtaion_2_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_2_booth_output_16, QB=>nx12676, D=>nx7091, CLK=>clk, 
      R=>rst);
   booth_integrtaion_2_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_2_15, QB=>nx12966, D=>nx7101, CLK=>clk, R=>
      rst);
   ix7887 : xor2 port map ( Y=>label_2(1), A0=>nx12983, A1=>nx12985);
   ix12984 : nand02 port map ( Y=>nx12983, A0=>adderInput_2(0), A1=>
      booth_integration_output_2_0);
   ix12986 : xnor2 port map ( Y=>nx12985, A0=>booth_integration_output_2_1, 
      A1=>adderInput_2(1));
   ix7885 : xor2 port map ( Y=>label_2(2), A0=>nx12988, A1=>nx12991);
   ix12989 : aoi32 port map ( Y=>nx12988, A0=>adderInput_2(0), A1=>
      booth_integration_output_2_0, A2=>nx7744, B0=>adderInput_2(1), B1=>
      booth_integration_output_2_1);
   ix7883 : xnor2 port map ( Y=>label_2(3), A0=>nx7758, A1=>nx12997);
   ix7759 : oai22 port map ( Y=>nx7758, A0=>nx12988, A1=>nx12991, B0=>
      nx12995, B1=>nx12980);
   ix12996 : inv01 port map ( Y=>nx12995, A=>adderInput_2(2));
   ix12998 : xnor2 port map ( Y=>nx12997, A0=>booth_integration_output_2_3, 
      A1=>adderInput_2(3));
   ix7881 : xor2 port map ( Y=>label_2(4), A0=>nx13000, A1=>nx13003);
   ix13001 : aoi22 port map ( Y=>nx13000, A0=>adderInput_2(3), A1=>
      booth_integration_output_2_3, B0=>nx7758, B1=>nx7760);
   ix7879 : xnor2 port map ( Y=>label_2(5), A0=>nx7774, A1=>nx13009);
   ix7775 : oai22 port map ( Y=>nx7774, A0=>nx13000, A1=>nx13003, B0=>
      nx13007, B1=>nx12978);
   ix13008 : inv01 port map ( Y=>nx13007, A=>adderInput_2(4));
   ix13010 : xnor2 port map ( Y=>nx13009, A0=>booth_integration_output_2_5, 
      A1=>adderInput_2(5));
   ix7877 : xor2 port map ( Y=>label_2(6), A0=>nx13012, A1=>nx13015);
   ix13013 : aoi22 port map ( Y=>nx13012, A0=>adderInput_2(5), A1=>
      booth_integration_output_2_5, B0=>nx7774, B1=>nx7776);
   ix7875 : xnor2 port map ( Y=>label_2(7), A0=>nx7790, A1=>nx13021);
   ix7791 : oai22 port map ( Y=>nx7790, A0=>nx13012, A1=>nx13015, B0=>
      nx13019, B1=>nx12976);
   ix13020 : inv01 port map ( Y=>nx13019, A=>adderInput_2(6));
   ix13022 : xnor2 port map ( Y=>nx13021, A0=>booth_integration_output_2_7, 
      A1=>adderInput_2(7));
   ix7873 : xor2 port map ( Y=>label_2(8), A0=>nx13024, A1=>nx13027);
   ix13025 : aoi22 port map ( Y=>nx13024, A0=>adderInput_2(7), A1=>
      booth_integration_output_2_7, B0=>nx7790, B1=>nx7792);
   ix7871 : xnor2 port map ( Y=>label_2(9), A0=>nx7806, A1=>nx13033);
   ix7807 : oai22 port map ( Y=>nx7806, A0=>nx13024, A1=>nx13027, B0=>
      nx13031, B1=>nx12974);
   ix13032 : inv01 port map ( Y=>nx13031, A=>adderInput_2(8));
   ix13034 : xnor2 port map ( Y=>nx13033, A0=>booth_integration_output_2_9, 
      A1=>adderInput_2(9));
   ix7869 : xor2 port map ( Y=>label_2(10), A0=>nx13036, A1=>nx13039);
   ix13037 : aoi22 port map ( Y=>nx13036, A0=>adderInput_2(9), A1=>
      booth_integration_output_2_9, B0=>nx7806, B1=>nx7808);
   ix7867 : xnor2 port map ( Y=>label_2(11), A0=>nx7822, A1=>nx13045);
   ix7823 : oai22 port map ( Y=>nx7822, A0=>nx13036, A1=>nx13039, B0=>
      nx13043, B1=>nx12972);
   ix13044 : inv01 port map ( Y=>nx13043, A=>adderInput_2(10));
   ix13046 : xnor2 port map ( Y=>nx13045, A0=>booth_integration_output_2_11, 
      A1=>adderInput_2(11));
   ix7865 : xor2 port map ( Y=>label_2(12), A0=>nx13048, A1=>nx13051);
   ix13049 : aoi22 port map ( Y=>nx13048, A0=>adderInput_2(11), A1=>
      booth_integration_output_2_11, B0=>nx7822, B1=>nx7824);
   ix7863 : xnor2 port map ( Y=>label_2(13), A0=>nx7838, A1=>nx13057);
   ix7839 : oai22 port map ( Y=>nx7838, A0=>nx13048, A1=>nx13051, B0=>
      nx13055, B1=>nx12970);
   ix13056 : inv01 port map ( Y=>nx13055, A=>adderInput_2(12));
   ix13058 : xnor2 port map ( Y=>nx13057, A0=>booth_integration_output_2_13, 
      A1=>adderInput_2(13));
   ix7861 : xor2 port map ( Y=>label_2(14), A0=>nx13060, A1=>nx13063);
   ix13061 : aoi22 port map ( Y=>nx13060, A0=>adderInput_2(13), A1=>
      booth_integration_output_2_13, B0=>nx7838, B1=>nx7840);
   ix7859 : xnor2 port map ( Y=>label_2(15), A0=>nx7854, A1=>nx13069);
   ix7855 : oai22 port map ( Y=>nx7854, A0=>nx13060, A1=>nx13063, B0=>
      nx13067, B1=>nx12968);
   ix13068 : inv01 port map ( Y=>nx13067, A=>adderInput_2(14));
   booth_integrtaion_1_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_1, QB=>OPEN, D=>nx7771, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_2, QB=>nx13503, D=>nx7761, CLK=>clk, R=>rst
   );
   booth_integrtaion_1_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_3, QB=>OPEN, D=>nx7751, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_4, QB=>nx13501, D=>nx7741, CLK=>clk, R=>rst
   );
   booth_integrtaion_1_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_5, QB=>OPEN, D=>nx7731, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_6, QB=>nx13499, D=>nx7721, CLK=>clk, R=>rst
   );
   booth_integrtaion_1_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_7, QB=>OPEN, D=>nx7711, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_8, QB=>nx13497, D=>nx7701, CLK=>clk, R=>rst
   );
   booth_integrtaion_1_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_9, QB=>OPEN, D=>nx7691, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_10, QB=>nx13495, D=>nx7681, CLK=>clk, R=>
      rst);
   booth_integrtaion_1_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_11, QB=>OPEN, D=>nx7671, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_12, QB=>nx13493, D=>nx7661, CLK=>clk, R=>
      rst);
   booth_integrtaion_1_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_13, QB=>OPEN, D=>nx7651, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_14, QB=>nx13491, D=>nx7641, CLK=>clk, R=>
      rst);
   ix13121 : aoi22 port map ( Y=>nx13120, A0=>neuron(15), A1=>nx14350, B0=>
      nx8530, B1=>nx8536);
   booth_integrtaion_1_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_reg_output_0, QB=>OPEN, D=>nx7281, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_0, QB=>OPEN, D=>nx7267, CLK=>clk, 
      S=>nx14168);
   booth_integrtaion_1_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_reg_output_9, QB=>OPEN, D=>nx7461, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_9, QB=>OPEN, D=>nx7451, CLK=>clk, 
      R=>nx14168);
   booth_integrtaion_1_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_8, QB=>OPEN, D=>nx7441, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_8, QB=>OPEN, D=>nx7431, CLK=>clk, 
      R=>nx14168);
   booth_integrtaion_1_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_7, QB=>OPEN, D=>nx7421, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_7, QB=>OPEN, D=>nx7411, CLK=>clk, 
      R=>nx14168);
   booth_integrtaion_1_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_6, QB=>OPEN, D=>nx7401, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_6, QB=>OPEN, D=>nx7391, CLK=>clk, 
      R=>nx14168);
   booth_integrtaion_1_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_5, QB=>OPEN, D=>nx7381, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_5, QB=>OPEN, D=>nx7371, CLK=>clk, 
      R=>nx14168);
   booth_integrtaion_1_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_4, QB=>OPEN, D=>nx7361, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_4, QB=>OPEN, D=>nx7351, CLK=>clk, 
      R=>nx14168);
   booth_integrtaion_1_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_3, QB=>OPEN, D=>nx7341, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_3, QB=>OPEN, D=>nx7331, CLK=>clk, 
      R=>nx14166);
   booth_integrtaion_1_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_2, QB=>OPEN, D=>nx7321, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_2, QB=>OPEN, D=>nx7311, CLK=>clk, 
      R=>nx14166);
   booth_integrtaion_1_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_output_1, QB=>OPEN, D=>nx7301, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_1_shift_Reg_count_1, QB=>OPEN, D=>nx7291, CLK=>clk, 
      R=>nx14166);
   ix7262 : nand02 port map ( Y=>nx7261, A0=>nx14644, A1=>nx14336);
   booth_integrtaion_1_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx13167, D=>nx7261, CLK=>clk, S=>nx14166);
   ix8531 : nand02 port map ( Y=>nx8530, A0=>nx13188, A1=>nx13199);
   ix13189 : oai21 port map ( Y=>nx13188, A0=>nx7994, A1=>nx7990, B0=>
      weight_1(0));
   ix7472 : oai21 port map ( Y=>nx7471, A0=>nx13193, A1=>nx14564, B0=>
      nx13195);
   booth_integrtaion_1_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13193, D=>nx7471, CLK=>clk, R=>rst);
   booth_integrtaion_1_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_0, QB=>nx13072, D=>nx7781, CLK=>clk, R=>rst
   );
   ix13204 : xnor2 port map ( Y=>nx13203, A0=>nx8000, A1=>nx2985);
   ix7612 : oai21 port map ( Y=>nx7611, A0=>nx13209, A1=>nx14564, B0=>
      nx13211);
   booth_integrtaion_1_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_17, QB=>nx13209, D=>nx7611, CLK=>clk, 
      R=>rst);
   ix13212 : nand03 port map ( Y=>nx13211, A0=>nx14572, A1=>nx8508, A2=>
      nx14786);
   ix8509 : xnor2 port map ( Y=>nx8508, A0=>nx13214, A1=>nx2986);
   ix13215 : aoi22 port map ( Y=>nx13214, A0=>
      booth_integrtaion_1_booth_output_17, A1=>nx8024, B0=>nx8000, B1=>
      nx2985);
   ix8009 : nand02 port map ( Y=>nx8008, A0=>weight_1(1), A1=>weight_1(0));
   ix13219 : or02 port map ( Y=>nx13218, A0=>weight_1(0), A1=>weight_1(1));
   ix7602 : oai21 port map ( Y=>nx7601, A0=>nx13223, A1=>nx14564, B0=>
      nx13225);
   booth_integrtaion_1_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13223, D=>nx7601, CLK=>clk, R=>rst);
   ix13226 : nand03 port map ( Y=>nx13225, A0=>nx14572, A1=>nx8496, A2=>
      nx14786);
   ix8497 : xnor2 port map ( Y=>nx8496, A0=>nx8052, A1=>nx13236);
   ix8053 : oai22 port map ( Y=>nx8052, A0=>nx13214, A1=>nx13229, B0=>
      nx13223, B1=>nx14576);
   ix13232 : aoi32 port map ( Y=>nx13231, A0=>nx8034, A1=>nx7994, A2=>
      nx13234, B0=>weight_1(2), B1=>nx7990);
   ix8035 : oai21 port map ( Y=>nx8034, A0=>weight_1(0), A1=>weight_1(1), B0
      =>weight_1(2));
   ix13237 : xnor2 port map ( Y=>nx13236, A0=>
      booth_integrtaion_1_booth_output_19, A1=>nx8072);
   booth_integrtaion_1_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_19, QB=>OPEN, D=>nx7591, CLK=>clk, R
      =>rst);
   ix13242 : xnor2 port map ( Y=>nx13241, A0=>nx13243, A1=>nx13257);
   ix13244 : aoi22 port map ( Y=>nx13243, A0=>
      booth_integrtaion_1_booth_output_19, A1=>nx8072, B0=>nx8052, B1=>
      nx2987);
   ix8073 : oai32 port map ( Y=>nx8072, A0=>nx13246, A1=>nx14578, A2=>nx8062, 
      B0=>nx13252, B1=>nx14582);
   ix13247 : nor02ii port map ( Y=>nx13246, A0=>nx8038, A1=>weight_1(3));
   ix8039 : nor03_2x port map ( Y=>nx8038, A0=>weight_1(2), A1=>weight_1(0), 
      A2=>weight_1(1));
   ix8063 : nor04 port map ( Y=>nx8062, A0=>weight_1(3), A1=>weight_1(2), A2
      =>weight_1(0), A3=>weight_1(1));
   ix13253 : inv01 port map ( Y=>nx13252, A=>weight_1(3));
   ix7582 : oai21 port map ( Y=>nx7581, A0=>nx13261, A1=>nx14564, B0=>
      nx13263);
   booth_integrtaion_1_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13261, D=>nx7581, CLK=>clk, R=>rst);
   ix13264 : nand03 port map ( Y=>nx13263, A0=>nx14572, A1=>nx8472, A2=>
      nx14786);
   ix8473 : xnor2 port map ( Y=>nx8472, A0=>nx8100, A1=>nx13276);
   ix8101 : oai22 port map ( Y=>nx8100, A0=>nx13243, A1=>nx13257, B0=>
      nx13261, B1=>nx13267);
   ix13275 : inv01 port map ( Y=>nx13274, A=>weight_1(4));
   ix13277 : xnor2 port map ( Y=>nx13276, A0=>
      booth_integrtaion_1_booth_output_21, A1=>nx8120);
   booth_integrtaion_1_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_21, QB=>OPEN, D=>nx7571, CLK=>clk, R
      =>rst);
   ix13282 : xnor2 port map ( Y=>nx13281, A0=>nx13283, A1=>nx13293);
   ix13284 : aoi22 port map ( Y=>nx13283, A0=>
      booth_integrtaion_1_booth_output_21, A1=>nx8120, B0=>nx8100, B1=>
      nx2989);
   ix8121 : oai32 port map ( Y=>nx8120, A0=>nx13286, A1=>nx14578, A2=>nx8110, 
      B0=>nx13290, B1=>nx14582);
   ix13287 : nor02ii port map ( Y=>nx13286, A0=>nx8086, A1=>weight_1(5));
   ix8087 : nor02ii port map ( Y=>nx8086, A0=>weight_1(4), A1=>nx8062);
   ix8111 : nor02ii port map ( Y=>nx8110, A0=>weight_1(5), A1=>nx8086);
   ix13291 : inv01 port map ( Y=>nx13290, A=>weight_1(5));
   ix7562 : oai21 port map ( Y=>nx7561, A0=>nx13297, A1=>nx14564, B0=>
      nx13299);
   booth_integrtaion_1_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13297, D=>nx7561, CLK=>clk, R=>rst);
   ix13300 : nand03 port map ( Y=>nx13299, A0=>nx14572, A1=>nx8448, A2=>
      nx14566);
   ix8449 : xnor2 port map ( Y=>nx8448, A0=>nx8148, A1=>nx13312);
   ix8149 : oai22 port map ( Y=>nx8148, A0=>nx13283, A1=>nx13293, B0=>
      nx13297, B1=>nx13303);
   ix13311 : inv01 port map ( Y=>nx13310, A=>weight_1(6));
   ix13313 : xnor2 port map ( Y=>nx13312, A0=>
      booth_integrtaion_1_booth_output_23, A1=>nx8168);
   booth_integrtaion_1_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_23, QB=>OPEN, D=>nx7551, CLK=>clk, R
      =>rst);
   ix13318 : xnor2 port map ( Y=>nx13317, A0=>nx13319, A1=>nx13329);
   ix13320 : aoi22 port map ( Y=>nx13319, A0=>
      booth_integrtaion_1_booth_output_23, A1=>nx8168, B0=>nx8148, B1=>
      nx2991);
   ix8169 : oai32 port map ( Y=>nx8168, A0=>nx13322, A1=>nx14578, A2=>nx8158, 
      B0=>nx13326, B1=>nx14582);
   ix13323 : nor02ii port map ( Y=>nx13322, A0=>nx8134, A1=>weight_1(7));
   ix8135 : nor02ii port map ( Y=>nx8134, A0=>weight_1(6), A1=>nx8110);
   ix8159 : nor02ii port map ( Y=>nx8158, A0=>weight_1(7), A1=>nx8134);
   ix13327 : inv01 port map ( Y=>nx13326, A=>weight_1(7));
   ix7542 : oai21 port map ( Y=>nx7541, A0=>nx13333, A1=>nx14566, B0=>
      nx13335);
   booth_integrtaion_1_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13333, D=>nx7541, CLK=>clk, R=>rst);
   ix13336 : nand03 port map ( Y=>nx13335, A0=>nx14572, A1=>nx8424, A2=>
      nx14566);
   ix8425 : xnor2 port map ( Y=>nx8424, A0=>nx8196, A1=>nx13348);
   ix8197 : oai22 port map ( Y=>nx8196, A0=>nx13319, A1=>nx13329, B0=>
      nx13333, B1=>nx13339);
   ix13347 : inv01 port map ( Y=>nx13346, A=>weight_1(8));
   ix13349 : xnor2 port map ( Y=>nx13348, A0=>
      booth_integrtaion_1_booth_output_25, A1=>nx8216);
   booth_integrtaion_1_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_25, QB=>OPEN, D=>nx7531, CLK=>clk, R
      =>rst);
   ix13354 : xnor2 port map ( Y=>nx13353, A0=>nx13355, A1=>nx13365);
   ix13356 : aoi22 port map ( Y=>nx13355, A0=>
      booth_integrtaion_1_booth_output_25, A1=>nx8216, B0=>nx8196, B1=>
      nx2993);
   ix8217 : oai32 port map ( Y=>nx8216, A0=>nx13358, A1=>nx14578, A2=>nx8206, 
      B0=>nx13362, B1=>nx14582);
   ix13359 : nor02ii port map ( Y=>nx13358, A0=>nx8182, A1=>weight_1(9));
   ix8183 : nor02ii port map ( Y=>nx8182, A0=>weight_1(8), A1=>nx8158);
   ix8207 : nor02ii port map ( Y=>nx8206, A0=>weight_1(9), A1=>nx8182);
   ix13363 : inv01 port map ( Y=>nx13362, A=>weight_1(9));
   ix7522 : oai21 port map ( Y=>nx7521, A0=>nx13369, A1=>nx14566, B0=>
      nx13371);
   booth_integrtaion_1_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13369, D=>nx7521, CLK=>clk, R=>rst);
   ix13372 : nand03 port map ( Y=>nx13371, A0=>nx14572, A1=>nx8400, A2=>
      nx14566);
   ix8401 : xnor2 port map ( Y=>nx8400, A0=>nx8244, A1=>nx13384);
   ix8245 : oai22 port map ( Y=>nx8244, A0=>nx13355, A1=>nx13365, B0=>
      nx13369, B1=>nx13375);
   ix13383 : inv01 port map ( Y=>nx13382, A=>weight_1(10));
   ix13385 : xnor2 port map ( Y=>nx13384, A0=>
      booth_integrtaion_1_booth_output_27, A1=>nx8264);
   booth_integrtaion_1_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_27, QB=>OPEN, D=>nx7511, CLK=>clk, R
      =>rst);
   ix13390 : xnor2 port map ( Y=>nx13389, A0=>nx13391, A1=>nx13401);
   ix13392 : aoi22 port map ( Y=>nx13391, A0=>
      booth_integrtaion_1_booth_output_27, A1=>nx8264, B0=>nx8244, B1=>
      nx2995);
   ix8265 : oai32 port map ( Y=>nx8264, A0=>nx13394, A1=>nx14578, A2=>nx8254, 
      B0=>nx13398, B1=>nx14582);
   ix13395 : nor02ii port map ( Y=>nx13394, A0=>nx8230, A1=>weight_1(11));
   ix8231 : nor02ii port map ( Y=>nx8230, A0=>weight_1(10), A1=>nx8206);
   ix8255 : nor02ii port map ( Y=>nx8254, A0=>weight_1(11), A1=>nx8230);
   ix13399 : inv01 port map ( Y=>nx13398, A=>weight_1(11));
   ix7502 : oai21 port map ( Y=>nx7501, A0=>nx13405, A1=>nx14566, B0=>
      nx13407);
   booth_integrtaion_1_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13405, D=>nx7501, CLK=>clk, R=>rst);
   ix13408 : nand03 port map ( Y=>nx13407, A0=>nx14794, A1=>nx8376, A2=>
      nx14566);
   ix8377 : xnor2 port map ( Y=>nx8376, A0=>nx8292, A1=>nx13420);
   ix8293 : oai22 port map ( Y=>nx8292, A0=>nx13391, A1=>nx13401, B0=>
      nx13405, B1=>nx13411);
   ix13419 : inv01 port map ( Y=>nx13418, A=>weight_1(12));
   ix13421 : xnor2 port map ( Y=>nx13420, A0=>
      booth_integrtaion_1_booth_output_29, A1=>nx8312);
   booth_integrtaion_1_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_29, QB=>OPEN, D=>nx7491, CLK=>clk, R
      =>rst);
   ix13426 : xnor2 port map ( Y=>nx13425, A0=>nx13427, A1=>nx13437);
   ix13428 : aoi22 port map ( Y=>nx13427, A0=>
      booth_integrtaion_1_booth_output_29, A1=>nx8312, B0=>nx8292, B1=>
      nx2997);
   ix8313 : oai32 port map ( Y=>nx8312, A0=>nx13430, A1=>nx14578, A2=>nx8302, 
      B0=>nx13434, B1=>nx14582);
   ix13431 : nor02ii port map ( Y=>nx13430, A0=>nx8278, A1=>weight_1(13));
   ix8279 : nor02ii port map ( Y=>nx8278, A0=>weight_1(12), A1=>nx8254);
   ix8303 : nor02ii port map ( Y=>nx8302, A0=>weight_1(13), A1=>nx8278);
   ix13435 : inv01 port map ( Y=>nx13434, A=>weight_1(13));
   ix13443 : xnor2 port map ( Y=>nx13442, A0=>nx8340, A1=>nx8350);
   ix8341 : oai22 port map ( Y=>nx8340, A0=>nx13427, A1=>nx13437, B0=>
      nx13445, B1=>nx13447);
   booth_integrtaion_1_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_31, QB=>nx13445, D=>nx7481, CLK=>clk, 
      R=>rst);
   ix13455 : inv01 port map ( Y=>nx13454, A=>weight_1(14));
   ix13458 : aoi22 port map ( Y=>nx13457, A0=>weight_1(15), A1=>nx7990, B0=>
      nx7994, B1=>nx8342);
   ix8343 : xnor2 port map ( Y=>nx8342, A0=>weight_1(15), A1=>nx8326);
   ix8327 : nor02ii port map ( Y=>nx8326, A0=>weight_1(14), A1=>nx8302);
   ix8337 : oai32 port map ( Y=>nx8336, A0=>nx13462, A1=>nx14578, A2=>nx8326, 
      B0=>nx13454, B1=>nx14582);
   ix13463 : nor02ii port map ( Y=>nx13462, A0=>nx8302, A1=>weight_1(14));
   ix8289 : oai32 port map ( Y=>nx8288, A0=>nx13466, A1=>nx14580, A2=>nx8278, 
      B0=>nx13418, B1=>nx14584);
   ix13467 : nor02ii port map ( Y=>nx13466, A0=>nx8254, A1=>weight_1(12));
   ix8241 : oai32 port map ( Y=>nx8240, A0=>nx13470, A1=>nx14580, A2=>nx8230, 
      B0=>nx13382, B1=>nx14584);
   ix13471 : nor02ii port map ( Y=>nx13470, A0=>nx8206, A1=>weight_1(10));
   ix8193 : oai32 port map ( Y=>nx8192, A0=>nx13474, A1=>nx14580, A2=>nx8182, 
      B0=>nx13346, B1=>nx14584);
   ix13475 : nor02ii port map ( Y=>nx13474, A0=>nx8158, A1=>weight_1(8));
   ix8145 : oai32 port map ( Y=>nx8144, A0=>nx13478, A1=>nx14580, A2=>nx8134, 
      B0=>nx13310, B1=>nx14584);
   ix13479 : nor02ii port map ( Y=>nx13478, A0=>nx8110, A1=>weight_1(6));
   ix8097 : oai32 port map ( Y=>nx8096, A0=>nx13482, A1=>nx14580, A2=>nx8086, 
      B0=>nx13274, B1=>nx14584);
   ix13483 : nor02ii port map ( Y=>nx13482, A0=>nx8062, A1=>weight_1(4));
   ix13486 : aoi32 port map ( Y=>nx13485, A0=>nx8008, A1=>nx7994, A2=>
      nx13218, B0=>weight_1(1), B1=>nx7990);
   booth_integrtaion_1_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_1_booth_output_16, QB=>nx13199, D=>nx7621, CLK=>clk, 
      R=>rst);
   booth_integrtaion_1_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_1_15, QB=>nx13489, D=>nx7631, CLK=>clk, R=>
      rst);
   ix8873 : xor2 port map ( Y=>label_1(1), A0=>nx13506, A1=>nx13508);
   ix13507 : nand02 port map ( Y=>nx13506, A0=>adderInput_1(0), A1=>
      booth_integration_output_1_0);
   ix13509 : xnor2 port map ( Y=>nx13508, A0=>booth_integration_output_1_1, 
      A1=>adderInput_1(1));
   ix8871 : xor2 port map ( Y=>label_1(2), A0=>nx13511, A1=>nx13514);
   ix13512 : aoi32 port map ( Y=>nx13511, A0=>adderInput_1(0), A1=>
      booth_integration_output_1_0, A2=>nx8730, B0=>adderInput_1(1), B1=>
      booth_integration_output_1_1);
   ix8869 : xnor2 port map ( Y=>label_1(3), A0=>nx8744, A1=>nx13520);
   ix8745 : oai22 port map ( Y=>nx8744, A0=>nx13511, A1=>nx13514, B0=>
      nx13518, B1=>nx13503);
   ix13519 : inv01 port map ( Y=>nx13518, A=>adderInput_1(2));
   ix13521 : xnor2 port map ( Y=>nx13520, A0=>booth_integration_output_1_3, 
      A1=>adderInput_1(3));
   ix8867 : xor2 port map ( Y=>label_1(4), A0=>nx13523, A1=>nx13526);
   ix13524 : aoi22 port map ( Y=>nx13523, A0=>adderInput_1(3), A1=>
      booth_integration_output_1_3, B0=>nx8744, B1=>nx8746);
   ix8865 : xnor2 port map ( Y=>label_1(5), A0=>nx8760, A1=>nx13532);
   ix8761 : oai22 port map ( Y=>nx8760, A0=>nx13523, A1=>nx13526, B0=>
      nx13530, B1=>nx13501);
   ix13531 : inv01 port map ( Y=>nx13530, A=>adderInput_1(4));
   ix13533 : xnor2 port map ( Y=>nx13532, A0=>booth_integration_output_1_5, 
      A1=>adderInput_1(5));
   ix8863 : xor2 port map ( Y=>label_1(6), A0=>nx13535, A1=>nx13538);
   ix13536 : aoi22 port map ( Y=>nx13535, A0=>adderInput_1(5), A1=>
      booth_integration_output_1_5, B0=>nx8760, B1=>nx8762);
   ix8861 : xnor2 port map ( Y=>label_1(7), A0=>nx8776, A1=>nx13544);
   ix8777 : oai22 port map ( Y=>nx8776, A0=>nx13535, A1=>nx13538, B0=>
      nx13542, B1=>nx13499);
   ix13543 : inv01 port map ( Y=>nx13542, A=>adderInput_1(6));
   ix13545 : xnor2 port map ( Y=>nx13544, A0=>booth_integration_output_1_7, 
      A1=>adderInput_1(7));
   ix8859 : xor2 port map ( Y=>label_1(8), A0=>nx13547, A1=>nx13550);
   ix13548 : aoi22 port map ( Y=>nx13547, A0=>adderInput_1(7), A1=>
      booth_integration_output_1_7, B0=>nx8776, B1=>nx8778);
   ix8857 : xnor2 port map ( Y=>label_1(9), A0=>nx8792, A1=>nx13556);
   ix8793 : oai22 port map ( Y=>nx8792, A0=>nx13547, A1=>nx13550, B0=>
      nx13554, B1=>nx13497);
   ix13555 : inv01 port map ( Y=>nx13554, A=>adderInput_1(8));
   ix13557 : xnor2 port map ( Y=>nx13556, A0=>booth_integration_output_1_9, 
      A1=>adderInput_1(9));
   ix8855 : xor2 port map ( Y=>label_1(10), A0=>nx13559, A1=>nx13562);
   ix13560 : aoi22 port map ( Y=>nx13559, A0=>adderInput_1(9), A1=>
      booth_integration_output_1_9, B0=>nx8792, B1=>nx8794);
   ix8853 : xnor2 port map ( Y=>label_1(11), A0=>nx8808, A1=>nx13568);
   ix8809 : oai22 port map ( Y=>nx8808, A0=>nx13559, A1=>nx13562, B0=>
      nx13566, B1=>nx13495);
   ix13567 : inv01 port map ( Y=>nx13566, A=>adderInput_1(10));
   ix13569 : xnor2 port map ( Y=>nx13568, A0=>booth_integration_output_1_11, 
      A1=>adderInput_1(11));
   ix8851 : xor2 port map ( Y=>label_1(12), A0=>nx13571, A1=>nx13574);
   ix13572 : aoi22 port map ( Y=>nx13571, A0=>adderInput_1(11), A1=>
      booth_integration_output_1_11, B0=>nx8808, B1=>nx8810);
   ix8849 : xnor2 port map ( Y=>label_1(13), A0=>nx8824, A1=>nx13580);
   ix8825 : oai22 port map ( Y=>nx8824, A0=>nx13571, A1=>nx13574, B0=>
      nx13578, B1=>nx13493);
   ix13579 : inv01 port map ( Y=>nx13578, A=>adderInput_1(12));
   ix13581 : xnor2 port map ( Y=>nx13580, A0=>booth_integration_output_1_13, 
      A1=>adderInput_1(13));
   ix8847 : xor2 port map ( Y=>label_1(14), A0=>nx13583, A1=>nx13586);
   ix13584 : aoi22 port map ( Y=>nx13583, A0=>adderInput_1(13), A1=>
      booth_integration_output_1_13, B0=>nx8824, B1=>nx8826);
   ix8845 : xnor2 port map ( Y=>label_1(15), A0=>nx8840, A1=>nx13592);
   ix8841 : oai22 port map ( Y=>nx8840, A0=>nx13583, A1=>nx13586, B0=>
      nx13590, B1=>nx13491);
   ix13591 : inv01 port map ( Y=>nx13590, A=>adderInput_1(14));
   booth_integrtaion_0_p_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_1, QB=>OPEN, D=>nx8301, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_2, QB=>nx14026, D=>nx8291, CLK=>clk, R=>rst
   );
   booth_integrtaion_0_p_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_3, QB=>OPEN, D=>nx8281, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_4, QB=>nx14024, D=>nx8271, CLK=>clk, R=>rst
   );
   booth_integrtaion_0_p_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_5, QB=>OPEN, D=>nx8261, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_6, QB=>nx14022, D=>nx8251, CLK=>clk, R=>rst
   );
   booth_integrtaion_0_p_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_7, QB=>OPEN, D=>nx8241, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_8, QB=>nx14020, D=>nx8231, CLK=>clk, R=>rst
   );
   booth_integrtaion_0_p_Reg_loop1_10_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_9, QB=>OPEN, D=>nx8221, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_11_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_10, QB=>nx14018, D=>nx8211, CLK=>clk, R=>
      rst);
   booth_integrtaion_0_p_Reg_loop1_12_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_11, QB=>OPEN, D=>nx8201, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_13_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_12, QB=>nx14016, D=>nx8191, CLK=>clk, R=>
      rst);
   booth_integrtaion_0_p_Reg_loop1_14_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_13, QB=>OPEN, D=>nx8181, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_15_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_14, QB=>nx14014, D=>nx8171, CLK=>clk, R=>
      rst);
   ix13644 : aoi22 port map ( Y=>nx13643, A0=>neuron(15), A1=>nx14372, B0=>
      nx9516, B1=>nx9522);
   booth_integrtaion_0_shift_Reg_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_reg_output_0, QB=>OPEN, D=>nx7811, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_0 : dffs_ni port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_0, QB=>OPEN, D=>nx7797, CLK=>clk, 
      S=>nx14172);
   booth_integrtaion_0_shift_Reg_Reg_loop1_9_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_reg_output_9, QB=>OPEN, D=>nx7991, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_9 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_9, QB=>OPEN, D=>nx7981, CLK=>clk, 
      R=>nx14172);
   booth_integrtaion_0_shift_Reg_Reg_loop1_8_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_8, QB=>OPEN, D=>nx7971, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_8 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_8, QB=>OPEN, D=>nx7961, CLK=>clk, 
      R=>nx14172);
   booth_integrtaion_0_shift_Reg_Reg_loop1_7_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_7, QB=>OPEN, D=>nx7951, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_7 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_7, QB=>OPEN, D=>nx7941, CLK=>clk, 
      R=>nx14172);
   booth_integrtaion_0_shift_Reg_Reg_loop1_6_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_6, QB=>OPEN, D=>nx7931, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_6 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_6, QB=>OPEN, D=>nx7921, CLK=>clk, 
      R=>nx14170);
   booth_integrtaion_0_shift_Reg_Reg_loop1_5_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_5, QB=>OPEN, D=>nx7911, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_5 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_5, QB=>OPEN, D=>nx7901, CLK=>clk, 
      R=>nx14170);
   booth_integrtaion_0_shift_Reg_Reg_loop1_4_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_4, QB=>OPEN, D=>nx7891, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_4 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_4, QB=>OPEN, D=>nx7881, CLK=>clk, 
      R=>nx14170);
   booth_integrtaion_0_shift_Reg_Reg_loop1_3_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_3, QB=>OPEN, D=>nx7871, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_3 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_3, QB=>OPEN, D=>nx7861, CLK=>clk, 
      R=>nx14170);
   booth_integrtaion_0_shift_Reg_Reg_loop1_2_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_2, QB=>OPEN, D=>nx7851, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_2 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_2, QB=>OPEN, D=>nx7841, CLK=>clk, 
      R=>nx14170);
   booth_integrtaion_0_shift_Reg_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_output_1, QB=>OPEN, D=>nx7831, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_shift_Reg_reg_count_1 : dffr port map ( Q=>
      booth_integrtaion_0_shift_Reg_count_1, QB=>OPEN, D=>nx7821, CLK=>clk, 
      R=>nx14170);
   ix7792 : nand02 port map ( Y=>nx7791, A0=>nx14648, A1=>nx14358);
   booth_integrtaion_0_shift_Reg_reg_en : dffs_ni port map ( Q=>OPEN, QB=>
      nx13690, D=>nx7791, CLK=>clk, S=>nx14170);
   ix9517 : nand02 port map ( Y=>nx9516, A0=>nx13711, A1=>nx13722);
   ix13712 : oai21 port map ( Y=>nx13711, A0=>nx8980, A1=>nx8976, B0=>
      weight_0(0));
   ix8002 : oai21 port map ( Y=>nx8001, A0=>nx13716, A1=>nx14586, B0=>
      nx13718);
   booth_integrtaion_0_p_Reg_loop1_0_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13716, D=>nx8001, CLK=>clk, R=>rst);
   booth_integrtaion_0_p_Reg_loop1_1_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_0, QB=>nx13595, D=>nx8311, CLK=>clk, R=>rst
   );
   ix13727 : xnor2 port map ( Y=>nx13726, A0=>nx8986, A1=>nx3000);
   ix8142 : oai21 port map ( Y=>nx8141, A0=>nx13732, A1=>nx14586, B0=>
      nx13734);
   booth_integrtaion_0_p_Reg_loop1_18_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_17, QB=>nx13732, D=>nx8141, CLK=>clk, 
      R=>rst);
   ix13735 : nand03 port map ( Y=>nx13734, A0=>nx14594, A1=>nx9494, A2=>
      nx14802);
   ix9495 : xnor2 port map ( Y=>nx9494, A0=>nx13737, A1=>nx3001);
   ix13738 : aoi22 port map ( Y=>nx13737, A0=>
      booth_integrtaion_0_booth_output_17, A1=>nx9010, B0=>nx8986, B1=>
      nx3000);
   ix8995 : nand02 port map ( Y=>nx8994, A0=>weight_0(1), A1=>weight_0(0));
   ix13742 : or02 port map ( Y=>nx13741, A0=>weight_0(0), A1=>weight_0(1));
   ix8132 : oai21 port map ( Y=>nx8131, A0=>nx13746, A1=>nx14586, B0=>
      nx13748);
   booth_integrtaion_0_p_Reg_loop1_19_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13746, D=>nx8131, CLK=>clk, R=>rst);
   ix13749 : nand03 port map ( Y=>nx13748, A0=>nx14594, A1=>nx9482, A2=>
      nx14802);
   ix9483 : xnor2 port map ( Y=>nx9482, A0=>nx9038, A1=>nx13759);
   ix9039 : oai22 port map ( Y=>nx9038, A0=>nx13737, A1=>nx13752, B0=>
      nx13746, B1=>nx14598);
   ix13755 : aoi32 port map ( Y=>nx13754, A0=>nx9020, A1=>nx8980, A2=>
      nx13757, B0=>weight_0(2), B1=>nx8976);
   ix9021 : oai21 port map ( Y=>nx9020, A0=>weight_0(0), A1=>weight_0(1), B0
      =>weight_0(2));
   ix13760 : xnor2 port map ( Y=>nx13759, A0=>
      booth_integrtaion_0_booth_output_19, A1=>nx9058);
   booth_integrtaion_0_p_Reg_loop1_20_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_19, QB=>OPEN, D=>nx8121, CLK=>clk, R
      =>rst);
   ix13765 : xnor2 port map ( Y=>nx13764, A0=>nx13766, A1=>nx13780);
   ix13767 : aoi22 port map ( Y=>nx13766, A0=>
      booth_integrtaion_0_booth_output_19, A1=>nx9058, B0=>nx9038, B1=>
      nx3002);
   ix9059 : oai32 port map ( Y=>nx9058, A0=>nx13769, A1=>nx14600, A2=>nx9048, 
      B0=>nx13775, B1=>nx14604);
   ix13770 : nor02ii port map ( Y=>nx13769, A0=>nx9024, A1=>weight_0(3));
   ix9025 : nor03_2x port map ( Y=>nx9024, A0=>weight_0(2), A1=>weight_0(0), 
      A2=>weight_0(1));
   ix9049 : nor04 port map ( Y=>nx9048, A0=>weight_0(3), A1=>weight_0(2), A2
      =>weight_0(0), A3=>weight_0(1));
   ix13776 : inv01 port map ( Y=>nx13775, A=>weight_0(3));
   ix8112 : oai21 port map ( Y=>nx8111, A0=>nx13784, A1=>nx14586, B0=>
      nx13786);
   booth_integrtaion_0_p_Reg_loop1_21_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13784, D=>nx8111, CLK=>clk, R=>rst);
   ix13787 : nand03 port map ( Y=>nx13786, A0=>nx14594, A1=>nx9458, A2=>
      nx14802);
   ix9459 : xnor2 port map ( Y=>nx9458, A0=>nx9086, A1=>nx13799);
   ix9087 : oai22 port map ( Y=>nx9086, A0=>nx13766, A1=>nx13780, B0=>
      nx13784, B1=>nx13790);
   ix13798 : inv01 port map ( Y=>nx13797, A=>weight_0(4));
   ix13800 : xnor2 port map ( Y=>nx13799, A0=>
      booth_integrtaion_0_booth_output_21, A1=>nx9106);
   booth_integrtaion_0_p_Reg_loop1_22_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_21, QB=>OPEN, D=>nx8101, CLK=>clk, R
      =>rst);
   ix13805 : xnor2 port map ( Y=>nx13804, A0=>nx13806, A1=>nx13816);
   ix13807 : aoi22 port map ( Y=>nx13806, A0=>
      booth_integrtaion_0_booth_output_21, A1=>nx9106, B0=>nx9086, B1=>
      nx3004);
   ix9107 : oai32 port map ( Y=>nx9106, A0=>nx13809, A1=>nx14600, A2=>nx9096, 
      B0=>nx13813, B1=>nx14604);
   ix13810 : nor02ii port map ( Y=>nx13809, A0=>nx9072, A1=>weight_0(5));
   ix9073 : nor02ii port map ( Y=>nx9072, A0=>weight_0(4), A1=>nx9048);
   ix9097 : nor02ii port map ( Y=>nx9096, A0=>weight_0(5), A1=>nx9072);
   ix13814 : inv01 port map ( Y=>nx13813, A=>weight_0(5));
   ix8092 : oai21 port map ( Y=>nx8091, A0=>nx13820, A1=>nx14586, B0=>
      nx13822);
   booth_integrtaion_0_p_Reg_loop1_23_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13820, D=>nx8091, CLK=>clk, R=>rst);
   ix13823 : nand03 port map ( Y=>nx13822, A0=>nx14594, A1=>nx9434, A2=>
      nx14588);
   ix9435 : xnor2 port map ( Y=>nx9434, A0=>nx9134, A1=>nx13835);
   ix9135 : oai22 port map ( Y=>nx9134, A0=>nx13806, A1=>nx13816, B0=>
      nx13820, B1=>nx13826);
   ix13834 : inv01 port map ( Y=>nx13833, A=>weight_0(6));
   ix13836 : xnor2 port map ( Y=>nx13835, A0=>
      booth_integrtaion_0_booth_output_23, A1=>nx9154);
   booth_integrtaion_0_p_Reg_loop1_24_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_23, QB=>OPEN, D=>nx8081, CLK=>clk, R
      =>rst);
   ix13841 : xnor2 port map ( Y=>nx13840, A0=>nx13842, A1=>nx13852);
   ix13843 : aoi22 port map ( Y=>nx13842, A0=>
      booth_integrtaion_0_booth_output_23, A1=>nx9154, B0=>nx9134, B1=>
      nx3006);
   ix9155 : oai32 port map ( Y=>nx9154, A0=>nx13845, A1=>nx14600, A2=>nx9144, 
      B0=>nx13849, B1=>nx14604);
   ix13846 : nor02ii port map ( Y=>nx13845, A0=>nx9120, A1=>weight_0(7));
   ix9121 : nor02ii port map ( Y=>nx9120, A0=>weight_0(6), A1=>nx9096);
   ix9145 : nor02ii port map ( Y=>nx9144, A0=>weight_0(7), A1=>nx9120);
   ix13850 : inv01 port map ( Y=>nx13849, A=>weight_0(7));
   ix8072 : oai21 port map ( Y=>nx8071, A0=>nx13856, A1=>nx14588, B0=>
      nx13858);
   booth_integrtaion_0_p_Reg_loop1_25_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13856, D=>nx8071, CLK=>clk, R=>rst);
   ix13859 : nand03 port map ( Y=>nx13858, A0=>nx14594, A1=>nx9410, A2=>
      nx14588);
   ix9411 : xnor2 port map ( Y=>nx9410, A0=>nx9182, A1=>nx13871);
   ix9183 : oai22 port map ( Y=>nx9182, A0=>nx13842, A1=>nx13852, B0=>
      nx13856, B1=>nx13862);
   ix13870 : inv01 port map ( Y=>nx13869, A=>weight_0(8));
   ix13872 : xnor2 port map ( Y=>nx13871, A0=>
      booth_integrtaion_0_booth_output_25, A1=>nx9202);
   booth_integrtaion_0_p_Reg_loop1_26_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_25, QB=>OPEN, D=>nx8061, CLK=>clk, R
      =>rst);
   ix13877 : xnor2 port map ( Y=>nx13876, A0=>nx13878, A1=>nx13888);
   ix13879 : aoi22 port map ( Y=>nx13878, A0=>
      booth_integrtaion_0_booth_output_25, A1=>nx9202, B0=>nx9182, B1=>
      nx3008);
   ix9203 : oai32 port map ( Y=>nx9202, A0=>nx13881, A1=>nx14600, A2=>nx9192, 
      B0=>nx13885, B1=>nx14604);
   ix13882 : nor02ii port map ( Y=>nx13881, A0=>nx9168, A1=>weight_0(9));
   ix9169 : nor02ii port map ( Y=>nx9168, A0=>weight_0(8), A1=>nx9144);
   ix9193 : nor02ii port map ( Y=>nx9192, A0=>weight_0(9), A1=>nx9168);
   ix13886 : inv01 port map ( Y=>nx13885, A=>weight_0(9));
   ix8052 : oai21 port map ( Y=>nx8051, A0=>nx13892, A1=>nx14588, B0=>
      nx13894);
   booth_integrtaion_0_p_Reg_loop1_27_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13892, D=>nx8051, CLK=>clk, R=>rst);
   ix13895 : nand03 port map ( Y=>nx13894, A0=>nx14594, A1=>nx9386, A2=>
      nx14588);
   ix9387 : xnor2 port map ( Y=>nx9386, A0=>nx9230, A1=>nx13907);
   ix9231 : oai22 port map ( Y=>nx9230, A0=>nx13878, A1=>nx13888, B0=>
      nx13892, B1=>nx13898);
   ix13906 : inv01 port map ( Y=>nx13905, A=>weight_0(10));
   ix13908 : xnor2 port map ( Y=>nx13907, A0=>
      booth_integrtaion_0_booth_output_27, A1=>nx9250);
   booth_integrtaion_0_p_Reg_loop1_28_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_27, QB=>OPEN, D=>nx8041, CLK=>clk, R
      =>rst);
   ix13913 : xnor2 port map ( Y=>nx13912, A0=>nx13914, A1=>nx13924);
   ix13915 : aoi22 port map ( Y=>nx13914, A0=>
      booth_integrtaion_0_booth_output_27, A1=>nx9250, B0=>nx9230, B1=>
      nx3010);
   ix9251 : oai32 port map ( Y=>nx9250, A0=>nx13917, A1=>nx14600, A2=>nx9240, 
      B0=>nx13921, B1=>nx14604);
   ix13918 : nor02ii port map ( Y=>nx13917, A0=>nx9216, A1=>weight_0(11));
   ix9217 : nor02ii port map ( Y=>nx9216, A0=>weight_0(10), A1=>nx9192);
   ix9241 : nor02ii port map ( Y=>nx9240, A0=>weight_0(11), A1=>nx9216);
   ix13922 : inv01 port map ( Y=>nx13921, A=>weight_0(11));
   ix8032 : oai21 port map ( Y=>nx8031, A0=>nx13928, A1=>nx14588, B0=>
      nx13930);
   booth_integrtaion_0_p_Reg_loop1_29_fx_reg_q : dffr port map ( Q=>OPEN, QB
      =>nx13928, D=>nx8031, CLK=>clk, R=>rst);
   ix13931 : nand03 port map ( Y=>nx13930, A0=>nx14810, A1=>nx9362, A2=>
      nx14588);
   ix9363 : xnor2 port map ( Y=>nx9362, A0=>nx9278, A1=>nx13943);
   ix9279 : oai22 port map ( Y=>nx9278, A0=>nx13914, A1=>nx13924, B0=>
      nx13928, B1=>nx13934);
   ix13942 : inv01 port map ( Y=>nx13941, A=>weight_0(12));
   ix13944 : xnor2 port map ( Y=>nx13943, A0=>
      booth_integrtaion_0_booth_output_29, A1=>nx9298);
   booth_integrtaion_0_p_Reg_loop1_30_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_29, QB=>OPEN, D=>nx8021, CLK=>clk, R
      =>rst);
   ix13949 : xnor2 port map ( Y=>nx13948, A0=>nx13950, A1=>nx13960);
   ix13951 : aoi22 port map ( Y=>nx13950, A0=>
      booth_integrtaion_0_booth_output_29, A1=>nx9298, B0=>nx9278, B1=>
      nx3012);
   ix9299 : oai32 port map ( Y=>nx9298, A0=>nx13953, A1=>nx14600, A2=>nx9288, 
      B0=>nx13957, B1=>nx14604);
   ix13954 : nor02ii port map ( Y=>nx13953, A0=>nx9264, A1=>weight_0(13));
   ix9265 : nor02ii port map ( Y=>nx9264, A0=>weight_0(12), A1=>nx9240);
   ix9289 : nor02ii port map ( Y=>nx9288, A0=>weight_0(13), A1=>nx9264);
   ix13958 : inv01 port map ( Y=>nx13957, A=>weight_0(13));
   ix13966 : xnor2 port map ( Y=>nx13965, A0=>nx9326, A1=>nx9336);
   ix9327 : oai22 port map ( Y=>nx9326, A0=>nx13950, A1=>nx13960, B0=>
      nx13968, B1=>nx13970);
   booth_integrtaion_0_p_Reg_loop1_32_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_31, QB=>nx13968, D=>nx8011, CLK=>clk, 
      R=>rst);
   ix13978 : inv01 port map ( Y=>nx13977, A=>weight_0(14));
   ix13981 : aoi22 port map ( Y=>nx13980, A0=>weight_0(15), A1=>nx8976, B0=>
      nx8980, B1=>nx9328);
   ix9329 : xnor2 port map ( Y=>nx9328, A0=>weight_0(15), A1=>nx9312);
   ix9313 : nor02ii port map ( Y=>nx9312, A0=>weight_0(14), A1=>nx9288);
   ix9323 : oai32 port map ( Y=>nx9322, A0=>nx13985, A1=>nx14600, A2=>nx9312, 
      B0=>nx13977, B1=>nx14604);
   ix13986 : nor02ii port map ( Y=>nx13985, A0=>nx9288, A1=>weight_0(14));
   ix9275 : oai32 port map ( Y=>nx9274, A0=>nx13989, A1=>nx14602, A2=>nx9264, 
      B0=>nx13941, B1=>nx14606);
   ix13990 : nor02ii port map ( Y=>nx13989, A0=>nx9240, A1=>weight_0(12));
   ix9227 : oai32 port map ( Y=>nx9226, A0=>nx13993, A1=>nx14602, A2=>nx9216, 
      B0=>nx13905, B1=>nx14606);
   ix13994 : nor02ii port map ( Y=>nx13993, A0=>nx9192, A1=>weight_0(10));
   ix9179 : oai32 port map ( Y=>nx9178, A0=>nx13997, A1=>nx14602, A2=>nx9168, 
      B0=>nx13869, B1=>nx14606);
   ix13998 : nor02ii port map ( Y=>nx13997, A0=>nx9144, A1=>weight_0(8));
   ix9131 : oai32 port map ( Y=>nx9130, A0=>nx14001, A1=>nx14602, A2=>nx9120, 
      B0=>nx13833, B1=>nx14606);
   ix14002 : nor02ii port map ( Y=>nx14001, A0=>nx9096, A1=>weight_0(6));
   ix9083 : oai32 port map ( Y=>nx9082, A0=>nx14005, A1=>nx14602, A2=>nx9072, 
      B0=>nx13797, B1=>nx14606);
   ix14006 : nor02ii port map ( Y=>nx14005, A0=>nx9048, A1=>weight_0(4));
   ix14009 : aoi32 port map ( Y=>nx14008, A0=>nx8994, A1=>nx8980, A2=>
      nx13741, B0=>weight_0(1), B1=>nx8976);
   booth_integrtaion_0_p_Reg_loop1_17_fx_reg_q : dffr port map ( Q=>
      booth_integrtaion_0_booth_output_16, QB=>nx13722, D=>nx8151, CLK=>clk, 
      R=>rst);
   booth_integrtaion_0_p_Reg_loop1_16_fx_reg_q : dffr port map ( Q=>
      booth_integration_output_0_15, QB=>nx14012, D=>nx8161, CLK=>clk, R=>
      rst);
   ix9859 : xor2 port map ( Y=>label_0(1), A0=>nx14029, A1=>nx14031);
   ix14030 : nand02 port map ( Y=>nx14029, A0=>adderInput_0(0), A1=>
      booth_integration_output_0_0);
   ix14032 : xnor2 port map ( Y=>nx14031, A0=>booth_integration_output_0_1, 
      A1=>adderInput_0(1));
   ix9857 : xor2 port map ( Y=>label_0(2), A0=>nx14034, A1=>nx14037);
   ix14035 : aoi32 port map ( Y=>nx14034, A0=>adderInput_0(0), A1=>
      booth_integration_output_0_0, A2=>nx9716, B0=>adderInput_0(1), B1=>
      booth_integration_output_0_1);
   ix9855 : xnor2 port map ( Y=>label_0(3), A0=>nx9730, A1=>nx14043);
   ix9731 : oai22 port map ( Y=>nx9730, A0=>nx14034, A1=>nx14037, B0=>
      nx14041, B1=>nx14026);
   ix14042 : inv01 port map ( Y=>nx14041, A=>adderInput_0(2));
   ix14044 : xnor2 port map ( Y=>nx14043, A0=>booth_integration_output_0_3, 
      A1=>adderInput_0(3));
   ix9853 : xor2 port map ( Y=>label_0(4), A0=>nx14046, A1=>nx14049);
   ix14047 : aoi22 port map ( Y=>nx14046, A0=>adderInput_0(3), A1=>
      booth_integration_output_0_3, B0=>nx9730, B1=>nx9732);
   ix9851 : xnor2 port map ( Y=>label_0(5), A0=>nx9746, A1=>nx14055);
   ix9747 : oai22 port map ( Y=>nx9746, A0=>nx14046, A1=>nx14049, B0=>
      nx14053, B1=>nx14024);
   ix14054 : inv01 port map ( Y=>nx14053, A=>adderInput_0(4));
   ix14056 : xnor2 port map ( Y=>nx14055, A0=>booth_integration_output_0_5, 
      A1=>adderInput_0(5));
   ix9849 : xor2 port map ( Y=>label_0(6), A0=>nx14058, A1=>nx14061);
   ix14059 : aoi22 port map ( Y=>nx14058, A0=>adderInput_0(5), A1=>
      booth_integration_output_0_5, B0=>nx9746, B1=>nx9748);
   ix9847 : xnor2 port map ( Y=>label_0(7), A0=>nx9762, A1=>nx14067);
   ix9763 : oai22 port map ( Y=>nx9762, A0=>nx14058, A1=>nx14061, B0=>
      nx14065, B1=>nx14022);
   ix14066 : inv01 port map ( Y=>nx14065, A=>adderInput_0(6));
   ix14068 : xnor2 port map ( Y=>nx14067, A0=>booth_integration_output_0_7, 
      A1=>adderInput_0(7));
   ix9845 : xor2 port map ( Y=>label_0(8), A0=>nx14070, A1=>nx14073);
   ix14071 : aoi22 port map ( Y=>nx14070, A0=>adderInput_0(7), A1=>
      booth_integration_output_0_7, B0=>nx9762, B1=>nx9764);
   ix9843 : xnor2 port map ( Y=>label_0(9), A0=>nx9778, A1=>nx14079);
   ix9779 : oai22 port map ( Y=>nx9778, A0=>nx14070, A1=>nx14073, B0=>
      nx14077, B1=>nx14020);
   ix14078 : inv01 port map ( Y=>nx14077, A=>adderInput_0(8));
   ix14080 : xnor2 port map ( Y=>nx14079, A0=>booth_integration_output_0_9, 
      A1=>adderInput_0(9));
   ix9841 : xor2 port map ( Y=>label_0(10), A0=>nx14082, A1=>nx14085);
   ix14083 : aoi22 port map ( Y=>nx14082, A0=>adderInput_0(9), A1=>
      booth_integration_output_0_9, B0=>nx9778, B1=>nx9780);
   ix9839 : xnor2 port map ( Y=>label_0(11), A0=>nx9794, A1=>nx14091);
   ix9795 : oai22 port map ( Y=>nx9794, A0=>nx14082, A1=>nx14085, B0=>
      nx14089, B1=>nx14018);
   ix14090 : inv01 port map ( Y=>nx14089, A=>adderInput_0(10));
   ix14092 : xnor2 port map ( Y=>nx14091, A0=>booth_integration_output_0_11, 
      A1=>adderInput_0(11));
   ix9837 : xor2 port map ( Y=>label_0(12), A0=>nx14094, A1=>nx14097);
   ix14095 : aoi22 port map ( Y=>nx14094, A0=>adderInput_0(11), A1=>
      booth_integration_output_0_11, B0=>nx9794, B1=>nx9796);
   ix9835 : xnor2 port map ( Y=>label_0(13), A0=>nx9810, A1=>nx14103);
   ix9811 : oai22 port map ( Y=>nx9810, A0=>nx14094, A1=>nx14097, B0=>
      nx14101, B1=>nx14016);
   ix14102 : inv01 port map ( Y=>nx14101, A=>adderInput_0(12));
   ix14104 : xnor2 port map ( Y=>nx14103, A0=>booth_integration_output_0_13, 
      A1=>adderInput_0(13));
   ix9833 : xor2 port map ( Y=>label_0(14), A0=>nx14106, A1=>nx14109);
   ix14107 : aoi22 port map ( Y=>nx14106, A0=>adderInput_0(13), A1=>
      booth_integration_output_0_13, B0=>nx9810, B1=>nx9812);
   ix9831 : xnor2 port map ( Y=>label_0(15), A0=>nx9826, A1=>nx14115);
   ix9827 : oai22 port map ( Y=>nx9826, A0=>nx14106, A1=>nx14109, B0=>
      nx14113, B1=>nx14014);
   ix14114 : inv01 port map ( Y=>nx14113, A=>adderInput_0(14));
   ix9813 : inv01 port map ( Y=>nx9812, A=>nx14103);
   ix9797 : inv01 port map ( Y=>nx9796, A=>nx14091);
   ix9781 : inv01 port map ( Y=>nx9780, A=>nx14079);
   ix9765 : inv01 port map ( Y=>nx9764, A=>nx14067);
   ix9749 : inv01 port map ( Y=>nx9748, A=>nx14055);
   ix9733 : inv01 port map ( Y=>nx9732, A=>nx14043);
   ix9717 : inv01 port map ( Y=>nx9716, A=>nx14031);
   ix13971 : inv01 port map ( Y=>nx13970, A=>nx9322);
   ix9361 : inv01 port map ( Y=>nx3012, A=>nx13943);
   ix13935 : inv01 port map ( Y=>nx13934, A=>nx9274);
   ix9385 : inv01 port map ( Y=>nx3010, A=>nx13907);
   ix13899 : inv01 port map ( Y=>nx13898, A=>nx9226);
   ix9409 : inv01 port map ( Y=>nx3008, A=>nx13871);
   ix13863 : inv01 port map ( Y=>nx13862, A=>nx9178);
   ix9433 : inv01 port map ( Y=>nx3006, A=>nx13835);
   ix13827 : inv01 port map ( Y=>nx13826, A=>nx9130);
   ix9457 : inv01 port map ( Y=>nx3004, A=>nx13799);
   ix13791 : inv01 port map ( Y=>nx13790, A=>nx9082);
   ix9481 : inv01 port map ( Y=>nx3002, A=>nx13759);
   ix13758 : inv01 port map ( Y=>nx13757, A=>nx9024);
   ix13753 : inv01 port map ( Y=>nx13752, A=>nx3001);
   ix9011 : inv01 port map ( Y=>nx9010, A=>nx14008);
   ix8827 : inv01 port map ( Y=>nx8826, A=>nx13580);
   ix8811 : inv01 port map ( Y=>nx8810, A=>nx13568);
   ix8795 : inv01 port map ( Y=>nx8794, A=>nx13556);
   ix8779 : inv01 port map ( Y=>nx8778, A=>nx13544);
   ix8763 : inv01 port map ( Y=>nx8762, A=>nx13532);
   ix8747 : inv01 port map ( Y=>nx8746, A=>nx13520);
   ix8731 : inv01 port map ( Y=>nx8730, A=>nx13508);
   ix13448 : inv01 port map ( Y=>nx13447, A=>nx8336);
   ix8375 : inv01 port map ( Y=>nx2997, A=>nx13420);
   ix13412 : inv01 port map ( Y=>nx13411, A=>nx8288);
   ix8399 : inv01 port map ( Y=>nx2995, A=>nx13384);
   ix13376 : inv01 port map ( Y=>nx13375, A=>nx8240);
   ix8423 : inv01 port map ( Y=>nx2993, A=>nx13348);
   ix13340 : inv01 port map ( Y=>nx13339, A=>nx8192);
   ix8447 : inv01 port map ( Y=>nx2991, A=>nx13312);
   ix13304 : inv01 port map ( Y=>nx13303, A=>nx8144);
   ix8471 : inv01 port map ( Y=>nx2989, A=>nx13276);
   ix13268 : inv01 port map ( Y=>nx13267, A=>nx8096);
   ix8495 : inv01 port map ( Y=>nx2987, A=>nx13236);
   ix13235 : inv01 port map ( Y=>nx13234, A=>nx8038);
   ix13230 : inv01 port map ( Y=>nx13229, A=>nx2986);
   ix8025 : inv01 port map ( Y=>nx8024, A=>nx13485);
   ix7841 : inv01 port map ( Y=>nx7840, A=>nx13057);
   ix7825 : inv01 port map ( Y=>nx7824, A=>nx13045);
   ix7809 : inv01 port map ( Y=>nx7808, A=>nx13033);
   ix7793 : inv01 port map ( Y=>nx7792, A=>nx13021);
   ix7777 : inv01 port map ( Y=>nx7776, A=>nx13009);
   ix7761 : inv01 port map ( Y=>nx7760, A=>nx12997);
   ix7745 : inv01 port map ( Y=>nx7744, A=>nx12985);
   ix12925 : inv01 port map ( Y=>nx12924, A=>nx7350);
   ix7389 : inv01 port map ( Y=>nx2982, A=>nx12897);
   ix12889 : inv01 port map ( Y=>nx12888, A=>nx7302);
   ix7413 : inv01 port map ( Y=>nx2980, A=>nx12861);
   ix12853 : inv01 port map ( Y=>nx12852, A=>nx7254);
   ix7437 : inv01 port map ( Y=>nx2978, A=>nx12825);
   ix12817 : inv01 port map ( Y=>nx12816, A=>nx7206);
   ix7461 : inv01 port map ( Y=>nx2976, A=>nx12789);
   ix12781 : inv01 port map ( Y=>nx12780, A=>nx7158);
   ix7485 : inv01 port map ( Y=>nx2974, A=>nx12753);
   ix12745 : inv01 port map ( Y=>nx12744, A=>nx7110);
   ix7509 : inv01 port map ( Y=>nx2972, A=>nx12713);
   ix12712 : inv01 port map ( Y=>nx12711, A=>nx7052);
   ix12707 : inv01 port map ( Y=>nx12706, A=>nx2971);
   ix7039 : inv01 port map ( Y=>nx7038, A=>nx12962);
   ix6855 : inv01 port map ( Y=>nx6854, A=>nx12534);
   ix6839 : inv01 port map ( Y=>nx6838, A=>nx12522);
   ix6823 : inv01 port map ( Y=>nx6822, A=>nx12510);
   ix6807 : inv01 port map ( Y=>nx6806, A=>nx12498);
   ix6791 : inv01 port map ( Y=>nx6790, A=>nx12486);
   ix6775 : inv01 port map ( Y=>nx6774, A=>nx12474);
   ix6759 : inv01 port map ( Y=>nx6758, A=>nx12462);
   ix12402 : inv01 port map ( Y=>nx12401, A=>nx6364);
   ix6403 : inv01 port map ( Y=>nx2967, A=>nx12374);
   ix12366 : inv01 port map ( Y=>nx12365, A=>nx6316);
   ix6427 : inv01 port map ( Y=>nx2965, A=>nx12338);
   ix12330 : inv01 port map ( Y=>nx12329, A=>nx6268);
   ix6451 : inv01 port map ( Y=>nx2963, A=>nx12302);
   ix12294 : inv01 port map ( Y=>nx12293, A=>nx6220);
   ix6475 : inv01 port map ( Y=>nx2961, A=>nx12266);
   ix12258 : inv01 port map ( Y=>nx12257, A=>nx6172);
   ix6499 : inv01 port map ( Y=>nx2959, A=>nx12230);
   ix12222 : inv01 port map ( Y=>nx12221, A=>nx6124);
   ix6523 : inv01 port map ( Y=>nx2956, A=>nx12190);
   ix12189 : inv01 port map ( Y=>nx12188, A=>nx6066);
   ix12184 : inv01 port map ( Y=>nx12183, A=>nx2955);
   ix6053 : inv01 port map ( Y=>nx6052, A=>nx12439);
   ix5869 : inv01 port map ( Y=>nx5868, A=>nx12011);
   ix5853 : inv01 port map ( Y=>nx5852, A=>nx11999);
   ix5837 : inv01 port map ( Y=>nx5836, A=>nx11987);
   ix5821 : inv01 port map ( Y=>nx5820, A=>nx11975);
   ix5805 : inv01 port map ( Y=>nx5804, A=>nx11963);
   ix5789 : inv01 port map ( Y=>nx5788, A=>nx11951);
   ix5773 : inv01 port map ( Y=>nx5772, A=>nx11939);
   ix11879 : inv01 port map ( Y=>nx11878, A=>nx5378);
   ix5417 : inv01 port map ( Y=>nx2951, A=>nx11851);
   ix11843 : inv01 port map ( Y=>nx11842, A=>nx5330);
   ix5441 : inv01 port map ( Y=>nx2949, A=>nx11815);
   ix11807 : inv01 port map ( Y=>nx11806, A=>nx5282);
   ix5465 : inv01 port map ( Y=>nx2947, A=>nx11779);
   ix11771 : inv01 port map ( Y=>nx11770, A=>nx5234);
   ix5489 : inv01 port map ( Y=>nx2945, A=>nx11743);
   ix11735 : inv01 port map ( Y=>nx11734, A=>nx5186);
   ix5513 : inv01 port map ( Y=>nx2943, A=>nx11707);
   ix11699 : inv01 port map ( Y=>nx11698, A=>nx5138);
   ix5537 : inv01 port map ( Y=>nx2941, A=>nx11667);
   ix11666 : inv01 port map ( Y=>nx11665, A=>nx5080);
   ix11661 : inv01 port map ( Y=>nx11660, A=>nx2940);
   ix5067 : inv01 port map ( Y=>nx5066, A=>nx11916);
   ix4883 : inv01 port map ( Y=>nx4882, A=>nx11488);
   ix4867 : inv01 port map ( Y=>nx4866, A=>nx11476);
   ix4851 : inv01 port map ( Y=>nx4850, A=>nx11464);
   ix4835 : inv01 port map ( Y=>nx4834, A=>nx11452);
   ix4819 : inv01 port map ( Y=>nx4818, A=>nx11440);
   ix4803 : inv01 port map ( Y=>nx4802, A=>nx11428);
   ix4787 : inv01 port map ( Y=>nx4786, A=>nx11416);
   ix11356 : inv01 port map ( Y=>nx11355, A=>nx4392);
   ix4431 : inv01 port map ( Y=>nx2936, A=>nx11328);
   ix11320 : inv01 port map ( Y=>nx11319, A=>nx4344);
   ix4455 : inv01 port map ( Y=>nx2934, A=>nx11292);
   ix11284 : inv01 port map ( Y=>nx11283, A=>nx4296);
   ix4479 : inv01 port map ( Y=>nx2932, A=>nx11256);
   ix11248 : inv01 port map ( Y=>nx11247, A=>nx4248);
   ix4503 : inv01 port map ( Y=>nx2930, A=>nx11220);
   ix11212 : inv01 port map ( Y=>nx11211, A=>nx4200);
   ix4527 : inv01 port map ( Y=>nx2928, A=>nx11184);
   ix11176 : inv01 port map ( Y=>nx11175, A=>nx4152);
   ix4551 : inv01 port map ( Y=>nx2925, A=>nx11144);
   ix11143 : inv01 port map ( Y=>nx11142, A=>nx4094);
   ix11138 : inv01 port map ( Y=>nx11137, A=>nx2923);
   ix4081 : inv01 port map ( Y=>nx4080, A=>nx11393);
   ix3897 : inv01 port map ( Y=>nx3896, A=>nx10965);
   ix3881 : inv01 port map ( Y=>nx3880, A=>nx10953);
   ix3865 : inv01 port map ( Y=>nx3864, A=>nx10941);
   ix3849 : inv01 port map ( Y=>nx3848, A=>nx10929);
   ix3833 : inv01 port map ( Y=>nx3832, A=>nx10917);
   ix3817 : inv01 port map ( Y=>nx3816, A=>nx10905);
   ix3801 : inv01 port map ( Y=>nx3800, A=>nx10893);
   ix10833 : inv01 port map ( Y=>nx10832, A=>nx3406);
   ix3445 : inv01 port map ( Y=>nx2915, A=>nx10805);
   ix10797 : inv01 port map ( Y=>nx10796, A=>nx3358);
   ix3469 : inv01 port map ( Y=>nx2911, A=>nx10769);
   ix10761 : inv01 port map ( Y=>nx10760, A=>nx3310);
   ix3493 : inv01 port map ( Y=>nx2907, A=>nx10733);
   ix10725 : inv01 port map ( Y=>nx10724, A=>nx3262);
   ix3517 : inv01 port map ( Y=>nx2903, A=>nx10697);
   ix10689 : inv01 port map ( Y=>nx10688, A=>nx3214);
   ix3541 : inv01 port map ( Y=>nx2899, A=>nx10661);
   ix10653 : inv01 port map ( Y=>nx10652, A=>nx3166);
   ix3565 : inv01 port map ( Y=>nx2895, A=>nx10621);
   ix10620 : inv01 port map ( Y=>nx10619, A=>nx3108);
   ix10615 : inv01 port map ( Y=>nx10614, A=>nx2893);
   ix3095 : inv01 port map ( Y=>nx3094, A=>nx10870);
   ix2911 : inv01 port map ( Y=>nx2910, A=>nx10442);
   ix2895 : inv01 port map ( Y=>nx2894, A=>nx10430);
   ix2879 : inv01 port map ( Y=>nx2878, A=>nx10418);
   ix2863 : inv01 port map ( Y=>nx2862, A=>nx10406);
   ix2847 : inv01 port map ( Y=>nx2846, A=>nx10394);
   ix2831 : inv01 port map ( Y=>nx2830, A=>nx10382);
   ix2815 : inv01 port map ( Y=>nx2814, A=>nx10370);
   ix10310 : inv01 port map ( Y=>nx10309, A=>nx2420);
   ix2459 : inv01 port map ( Y=>nx2885, A=>nx10282);
   ix10274 : inv01 port map ( Y=>nx10273, A=>nx2372);
   ix2483 : inv01 port map ( Y=>nx2881, A=>nx10246);
   ix10238 : inv01 port map ( Y=>nx10237, A=>nx2324);
   ix2507 : inv01 port map ( Y=>nx2877, A=>nx10210);
   ix10202 : inv01 port map ( Y=>nx10201, A=>nx2276);
   ix2531 : inv01 port map ( Y=>nx2873, A=>nx10174);
   ix10166 : inv01 port map ( Y=>nx10165, A=>nx2228);
   ix2555 : inv01 port map ( Y=>nx2869, A=>nx10138);
   ix10130 : inv01 port map ( Y=>nx10129, A=>nx2180);
   ix2579 : inv01 port map ( Y=>nx2865, A=>nx10098);
   ix10097 : inv01 port map ( Y=>nx10096, A=>nx2122);
   ix10092 : inv01 port map ( Y=>nx10091, A=>nx2863);
   ix2109 : inv01 port map ( Y=>nx2108, A=>nx10347);
   ix1925 : inv01 port map ( Y=>nx1924, A=>nx9919);
   ix1909 : inv01 port map ( Y=>nx1908, A=>nx9907);
   ix1893 : inv01 port map ( Y=>nx1892, A=>nx9895);
   ix1877 : inv01 port map ( Y=>nx1876, A=>nx9883);
   ix1861 : inv01 port map ( Y=>nx1860, A=>nx9870);
   ix1845 : inv01 port map ( Y=>nx1844, A=>nx9855);
   ix1829 : inv01 port map ( Y=>nx1828, A=>nx9839);
   ix9762 : inv01 port map ( Y=>nx9761, A=>nx1434);
   ix1473 : inv01 port map ( Y=>nx2855, A=>nx9723);
   ix9714 : inv01 port map ( Y=>nx9713, A=>nx1386);
   ix1497 : inv01 port map ( Y=>nx2851, A=>nx9681);
   ix9672 : inv01 port map ( Y=>nx9671, A=>nx1338);
   ix1521 : inv01 port map ( Y=>nx2847, A=>nx9639);
   ix9630 : inv01 port map ( Y=>nx9629, A=>nx1290);
   ix1545 : inv01 port map ( Y=>nx2843, A=>nx9595);
   ix9586 : inv01 port map ( Y=>nx9585, A=>nx1242);
   ix1569 : inv01 port map ( Y=>nx2839, A=>nx9553);
   ix9545 : inv01 port map ( Y=>nx9544, A=>nx1194);
   ix1593 : inv01 port map ( Y=>nx2835, A=>nx9507);
   ix9506 : inv01 port map ( Y=>nx9504, A=>nx1136);
   ix9500 : inv01 port map ( Y=>nx9499, A=>nx2833);
   ix1123 : inv01 port map ( Y=>nx1122, A=>nx9805);
   ix939 : inv01 port map ( Y=>nx938, A=>nx9263);
   ix923 : inv01 port map ( Y=>nx922, A=>nx9247);
   ix907 : inv01 port map ( Y=>nx906, A=>nx9231);
   ix891 : inv01 port map ( Y=>nx890, A=>nx9215);
   ix875 : inv01 port map ( Y=>nx874, A=>nx9199);
   ix859 : inv01 port map ( Y=>nx858, A=>nx9183);
   ix843 : inv01 port map ( Y=>nx842, A=>nx9167);
   ix9090 : inv01 port map ( Y=>nx9089, A=>nx448);
   ix487 : inv01 port map ( Y=>nx2825, A=>nx9051);
   ix9042 : inv01 port map ( Y=>nx9041, A=>nx400);
   ix511 : inv01 port map ( Y=>nx2821, A=>nx9003);
   ix8994 : inv01 port map ( Y=>nx8993, A=>nx352);
   ix535 : inv01 port map ( Y=>nx2817, A=>nx8960);
   ix8952 : inv01 port map ( Y=>nx8951, A=>nx304);
   ix559 : inv01 port map ( Y=>nx2813, A=>nx8924);
   ix8916 : inv01 port map ( Y=>nx8915, A=>nx256);
   ix583 : inv01 port map ( Y=>nx2810, A=>nx8888);
   ix8880 : inv01 port map ( Y=>nx8879, A=>nx208);
   ix607 : inv01 port map ( Y=>nx2808, A=>nx8837);
   ix8836 : inv01 port map ( Y=>nx8835, A=>nx150);
   ix8830 : inv01 port map ( Y=>nx8829, A=>nx2807);
   ix137 : inv01 port map ( Y=>nx136, A=>nx9133);
   ix14121 : inv02 port map ( Y=>nx14122, A=>nx14658);
   ix14135 : inv02 port map ( Y=>nx14136, A=>set);
   ix14137 : inv02 port map ( Y=>nx14138, A=>set);
   ix14139 : inv02 port map ( Y=>nx14140, A=>set);
   ix14141 : inv02 port map ( Y=>nx14142, A=>set);
   ix14143 : inv02 port map ( Y=>nx14144, A=>set);
   ix14145 : inv02 port map ( Y=>nx14146, A=>set);
   ix14147 : inv02 port map ( Y=>nx14148, A=>set);
   ix14149 : inv02 port map ( Y=>nx14150, A=>set);
   ix14151 : inv02 port map ( Y=>nx14152, A=>set);
   ix14153 : inv02 port map ( Y=>nx14154, A=>set);
   ix14155 : inv02 port map ( Y=>nx14156, A=>set);
   ix14157 : inv02 port map ( Y=>nx14158, A=>set);
   ix14159 : inv02 port map ( Y=>nx14160, A=>set);
   ix14161 : inv02 port map ( Y=>nx14162, A=>set);
   ix14163 : inv02 port map ( Y=>nx14164, A=>set);
   ix14165 : inv02 port map ( Y=>nx14166, A=>set);
   ix14167 : inv02 port map ( Y=>nx14168, A=>set);
   ix14169 : inv02 port map ( Y=>nx14170, A=>set);
   ix14171 : inv02 port map ( Y=>nx14172, A=>set);
   ix14173 : inv02 port map ( Y=>nx14174, A=>nx14666);
   ix14181 : inv02 port map ( Y=>nx14182, A=>nx14674);
   ix14195 : inv02 port map ( Y=>nx14196, A=>nx14682);
   ix14203 : inv02 port map ( Y=>nx14204, A=>nx14690);
   ix14217 : inv02 port map ( Y=>nx14218, A=>nx14698);
   ix14225 : inv02 port map ( Y=>nx14226, A=>nx14706);
   ix14239 : inv02 port map ( Y=>nx14240, A=>nx14714);
   ix14247 : inv02 port map ( Y=>nx14248, A=>nx14722);
   ix14261 : inv02 port map ( Y=>nx14262, A=>nx14730);
   ix14269 : inv02 port map ( Y=>nx14270, A=>nx14738);
   ix14283 : inv02 port map ( Y=>nx14284, A=>nx14746);
   ix14291 : inv02 port map ( Y=>nx14292, A=>nx14754);
   ix14305 : inv02 port map ( Y=>nx14306, A=>nx14762);
   ix14313 : inv02 port map ( Y=>nx14314, A=>nx14770);
   ix14327 : inv02 port map ( Y=>nx14328, A=>nx14778);
   ix14335 : inv02 port map ( Y=>nx14336, A=>nx14786);
   ix14349 : inv02 port map ( Y=>nx14350, A=>nx14794);
   ix14357 : inv02 port map ( Y=>nx14358, A=>nx14802);
   ix14371 : inv02 port map ( Y=>nx14372, A=>nx14810);
   ix14381 : inv02 port map ( Y=>nx14382, A=>nx14652);
   ix14387 : inv02 port map ( Y=>nx14388, A=>
      booth_integrtaion_9_shift_reg_output_9);
   ix14389 : inv02 port map ( Y=>nx14390, A=>nx14822);
   ix14391 : inv02 port map ( Y=>nx14392, A=>nx14822);
   ix14393 : inv02 port map ( Y=>nx14394, A=>nx14822);
   ix14395 : inv01 port map ( Y=>nx14396, A=>
      booth_integrtaion_9_shift_reg_output_0);
   ix14399 : buf02 port map ( Y=>nx14400, A=>nx8831);
   ix14401 : inv02 port map ( Y=>nx14402, A=>nx106);
   ix14403 : inv02 port map ( Y=>nx14404, A=>nx106);
   ix14405 : inv02 port map ( Y=>nx14406, A=>nx102);
   ix14407 : inv02 port map ( Y=>nx14408, A=>nx102);
   ix14409 : inv02 port map ( Y=>nx14410, A=>
      booth_integrtaion_8_shift_reg_output_9);
   ix14411 : inv02 port map ( Y=>nx14412, A=>nx14826);
   ix14413 : inv02 port map ( Y=>nx14414, A=>nx14826);
   ix14415 : inv02 port map ( Y=>nx14416, A=>nx14826);
   ix14417 : inv01 port map ( Y=>nx14418, A=>
      booth_integrtaion_8_shift_reg_output_0);
   ix14421 : buf02 port map ( Y=>nx14422, A=>nx9501);
   ix14423 : inv02 port map ( Y=>nx14424, A=>nx1092);
   ix14425 : inv02 port map ( Y=>nx14426, A=>nx1092);
   ix14427 : inv02 port map ( Y=>nx14428, A=>nx1088);
   ix14429 : inv02 port map ( Y=>nx14430, A=>nx1088);
   ix14431 : inv02 port map ( Y=>nx14432, A=>
      booth_integrtaion_7_shift_reg_output_9);
   ix14433 : inv02 port map ( Y=>nx14434, A=>nx14830);
   ix14435 : inv02 port map ( Y=>nx14436, A=>nx14830);
   ix14437 : inv02 port map ( Y=>nx14438, A=>nx14830);
   ix14439 : inv01 port map ( Y=>nx14440, A=>
      booth_integrtaion_7_shift_reg_output_0);
   ix14443 : buf02 port map ( Y=>nx14444, A=>nx10093);
   ix14445 : inv02 port map ( Y=>nx14446, A=>nx2078);
   ix14447 : inv02 port map ( Y=>nx14448, A=>nx2078);
   ix14449 : inv02 port map ( Y=>nx14450, A=>nx2074);
   ix14451 : inv02 port map ( Y=>nx14452, A=>nx2074);
   ix14453 : inv02 port map ( Y=>nx14454, A=>
      booth_integrtaion_6_shift_reg_output_9);
   ix14455 : inv02 port map ( Y=>nx14456, A=>nx14834);
   ix14457 : inv02 port map ( Y=>nx14458, A=>nx14834);
   ix14459 : inv02 port map ( Y=>nx14460, A=>nx14834);
   ix14461 : inv01 port map ( Y=>nx14462, A=>
      booth_integrtaion_6_shift_reg_output_0);
   ix14465 : buf02 port map ( Y=>nx14466, A=>nx10616);
   ix14467 : inv02 port map ( Y=>nx14468, A=>nx3064);
   ix14469 : inv02 port map ( Y=>nx14470, A=>nx3064);
   ix14471 : inv02 port map ( Y=>nx14472, A=>nx3060);
   ix14473 : inv02 port map ( Y=>nx14474, A=>nx3060);
   ix14475 : inv02 port map ( Y=>nx14476, A=>
      booth_integrtaion_5_shift_reg_output_9);
   ix14477 : inv02 port map ( Y=>nx14478, A=>nx14838);
   ix14479 : inv02 port map ( Y=>nx14480, A=>nx14838);
   ix14481 : inv02 port map ( Y=>nx14482, A=>nx14838);
   ix14483 : inv01 port map ( Y=>nx14484, A=>
      booth_integrtaion_5_shift_reg_output_0);
   ix14487 : buf02 port map ( Y=>nx14488, A=>nx11139);
   ix14489 : inv02 port map ( Y=>nx14490, A=>nx4050);
   ix14491 : inv02 port map ( Y=>nx14492, A=>nx4050);
   ix14493 : inv02 port map ( Y=>nx14494, A=>nx4046);
   ix14495 : inv02 port map ( Y=>nx14496, A=>nx4046);
   ix14497 : inv02 port map ( Y=>nx14498, A=>
      booth_integrtaion_4_shift_reg_output_9);
   ix14499 : inv02 port map ( Y=>nx14500, A=>nx14842);
   ix14501 : inv02 port map ( Y=>nx14502, A=>nx14842);
   ix14503 : inv02 port map ( Y=>nx14504, A=>nx14842);
   ix14505 : inv01 port map ( Y=>nx14506, A=>
      booth_integrtaion_4_shift_reg_output_0);
   ix14509 : buf02 port map ( Y=>nx14510, A=>nx11662);
   ix14511 : inv02 port map ( Y=>nx14512, A=>nx5036);
   ix14513 : inv02 port map ( Y=>nx14514, A=>nx5036);
   ix14515 : inv02 port map ( Y=>nx14516, A=>nx5032);
   ix14517 : inv02 port map ( Y=>nx14518, A=>nx5032);
   ix14519 : inv02 port map ( Y=>nx14520, A=>
      booth_integrtaion_3_shift_reg_output_9);
   ix14521 : inv02 port map ( Y=>nx14522, A=>nx14846);
   ix14523 : inv02 port map ( Y=>nx14524, A=>nx14846);
   ix14525 : inv02 port map ( Y=>nx14526, A=>nx14846);
   ix14527 : inv01 port map ( Y=>nx14528, A=>
      booth_integrtaion_3_shift_reg_output_0);
   ix14531 : buf02 port map ( Y=>nx14532, A=>nx12185);
   ix14533 : inv02 port map ( Y=>nx14534, A=>nx6022);
   ix14535 : inv02 port map ( Y=>nx14536, A=>nx6022);
   ix14537 : inv02 port map ( Y=>nx14538, A=>nx6018);
   ix14539 : inv02 port map ( Y=>nx14540, A=>nx6018);
   ix14541 : inv02 port map ( Y=>nx14542, A=>
      booth_integrtaion_2_shift_reg_output_9);
   ix14543 : inv02 port map ( Y=>nx14544, A=>nx14850);
   ix14545 : inv02 port map ( Y=>nx14546, A=>nx14850);
   ix14547 : inv02 port map ( Y=>nx14548, A=>nx14850);
   ix14549 : inv01 port map ( Y=>nx14550, A=>
      booth_integrtaion_2_shift_reg_output_0);
   ix14553 : buf02 port map ( Y=>nx14554, A=>nx12708);
   ix14555 : inv02 port map ( Y=>nx14556, A=>nx7008);
   ix14557 : inv02 port map ( Y=>nx14558, A=>nx7008);
   ix14559 : inv02 port map ( Y=>nx14560, A=>nx7004);
   ix14561 : inv02 port map ( Y=>nx14562, A=>nx7004);
   ix14563 : inv02 port map ( Y=>nx14564, A=>
      booth_integrtaion_1_shift_reg_output_9);
   ix14565 : inv02 port map ( Y=>nx14566, A=>nx14854);
   ix14567 : inv02 port map ( Y=>nx14568, A=>nx14854);
   ix14569 : inv02 port map ( Y=>nx14570, A=>nx14854);
   ix14571 : inv01 port map ( Y=>nx14572, A=>
      booth_integrtaion_1_shift_reg_output_0);
   ix14575 : buf02 port map ( Y=>nx14576, A=>nx13231);
   ix14577 : inv02 port map ( Y=>nx14578, A=>nx7994);
   ix14579 : inv02 port map ( Y=>nx14580, A=>nx7994);
   ix14581 : inv02 port map ( Y=>nx14582, A=>nx7990);
   ix14583 : inv02 port map ( Y=>nx14584, A=>nx7990);
   ix14585 : inv02 port map ( Y=>nx14586, A=>
      booth_integrtaion_0_shift_reg_output_9);
   ix14587 : inv02 port map ( Y=>nx14588, A=>nx14858);
   ix14589 : inv02 port map ( Y=>nx14590, A=>nx14858);
   ix14591 : inv02 port map ( Y=>nx14592, A=>nx14858);
   ix14593 : inv01 port map ( Y=>nx14594, A=>
      booth_integrtaion_0_shift_reg_output_0);
   ix14597 : buf02 port map ( Y=>nx14598, A=>nx13754);
   ix14599 : inv02 port map ( Y=>nx14600, A=>nx8980);
   ix14601 : inv02 port map ( Y=>nx14602, A=>nx8980);
   ix14603 : inv02 port map ( Y=>nx14604, A=>nx8976);
   ix14605 : inv02 port map ( Y=>nx14606, A=>nx8976);
   ix8512 : mux21_ni port map ( Y=>nx8511, A0=>dec_sel_0_EXMPLR, A1=>
      shift_Reg_adder_0_output_17, S0=>nx14652);
   ix8502 : mux21_ni port map ( Y=>nx8501, A0=>shift_Reg_adder_0_output_17, 
      A1=>shift_Reg_adder_0_output_16, S0=>nx14652);
   ix8492 : mux21_ni port map ( Y=>nx8491, A0=>shift_Reg_adder_0_output_16, 
      A1=>shift_Reg_adder_0_output_15, S0=>nx14652);
   ix8482 : mux21_ni port map ( Y=>nx8481, A0=>shift_Reg_adder_0_output_15, 
      A1=>shift_Reg_adder_0_output_14, S0=>nx14652);
   ix8472 : mux21_ni port map ( Y=>nx8471, A0=>shift_Reg_adder_0_output_14, 
      A1=>shift_Reg_adder_0_output_13, S0=>nx14652);
   ix8462 : mux21_ni port map ( Y=>nx8461, A0=>shift_Reg_adder_0_output_13, 
      A1=>shift_Reg_adder_0_output_12, S0=>nx14652);
   ix8452 : mux21_ni port map ( Y=>nx8451, A0=>shift_Reg_adder_0_output_12, 
      A1=>shift_Reg_adder_0_output_11, S0=>nx14654);
   ix8442 : mux21_ni port map ( Y=>nx8441, A0=>shift_Reg_adder_0_output_11, 
      A1=>shift_Reg_adder_0_output_10, S0=>nx14654);
   ix8432 : mux21_ni port map ( Y=>nx8431, A0=>shift_Reg_adder_0_output_10, 
      A1=>shift_Reg_adder_0_output_9, S0=>nx14654);
   ix8422 : mux21_ni port map ( Y=>nx8421, A0=>shift_Reg_adder_0_output_9, 
      A1=>shift_Reg_adder_0_output_8, S0=>nx14654);
   ix8412 : mux21_ni port map ( Y=>nx8411, A0=>shift_Reg_adder_0_output_8, 
      A1=>shift_Reg_adder_0_output_7, S0=>nx14654);
   ix8402 : mux21_ni port map ( Y=>nx8401, A0=>shift_Reg_adder_0_output_7, 
      A1=>shift_Reg_adder_0_output_6, S0=>nx14654);
   ix8392 : mux21_ni port map ( Y=>nx8391, A0=>shift_Reg_adder_0_output_6, 
      A1=>shift_Reg_adder_0_output_5, S0=>nx14654);
   ix8382 : mux21_ni port map ( Y=>nx8381, A0=>shift_Reg_adder_0_output_5, 
      A1=>shift_Reg_adder_0_output_4, S0=>nx14656);
   ix8372 : mux21_ni port map ( Y=>nx8371, A0=>shift_Reg_adder_0_output_4, 
      A1=>shift_Reg_adder_0_output_3, S0=>nx14656);
   ix8362 : mux21_ni port map ( Y=>nx8361, A0=>shift_Reg_adder_0_output_3, 
      A1=>shift_Reg_adder_0_output_2, S0=>nx14656);
   ix8352 : mux21_ni port map ( Y=>nx8351, A0=>shift_Reg_adder_0_output_2, 
      A1=>shift_Reg_adder_0_output_1, S0=>nx14656);
   ix8342 : mux21_ni port map ( Y=>nx8341, A0=>shift_Reg_adder_0_output_1, 
      A1=>shift_Reg_adder_0_output_0, S0=>nx14656);
   ix8328 : nor02ii port map ( Y=>nx8327, A0=>nx14656, A1=>
      shift_Reg_adder_0_output_0);
   ix991 : xor2 port map ( Y=>label_9(0), A0=>adderInput_9(0), A1=>
      booth_integration_output_9_0);
   ix3542 : mux21_ni port map ( Y=>nx3541, A0=>booth_integration_output_9_0, 
      A1=>nx834, S0=>nx14394);
   ix835 : mux21_ni port map ( Y=>nx834, A0=>neuron(0), A1=>
      booth_integration_output_9_1, S0=>nx14666);
   ix3532 : mux21_ni port map ( Y=>nx3531, A0=>booth_integration_output_9_1, 
      A1=>nx822, S0=>nx14394);
   ix823 : mux21_ni port map ( Y=>nx822, A0=>neuron(1), A1=>
      booth_integration_output_9_2, S0=>nx14666);
   ix3522 : mux21_ni port map ( Y=>nx3521, A0=>booth_integration_output_9_2, 
      A1=>nx810, S0=>nx14394);
   ix811 : mux21_ni port map ( Y=>nx810, A0=>neuron(2), A1=>
      booth_integration_output_9_3, S0=>nx14666);
   ix3512 : mux21_ni port map ( Y=>nx3511, A0=>booth_integration_output_9_3, 
      A1=>nx798, S0=>nx14394);
   ix799 : mux21_ni port map ( Y=>nx798, A0=>neuron(3), A1=>
      booth_integration_output_9_4, S0=>nx14666);
   ix3502 : mux21_ni port map ( Y=>nx3501, A0=>booth_integration_output_9_4, 
      A1=>nx786, S0=>nx14394);
   ix787 : mux21_ni port map ( Y=>nx786, A0=>neuron(4), A1=>
      booth_integration_output_9_5, S0=>nx14666);
   ix3492 : mux21_ni port map ( Y=>nx3491, A0=>booth_integration_output_9_5, 
      A1=>nx774, S0=>nx14394);
   ix775 : mux21_ni port map ( Y=>nx774, A0=>neuron(5), A1=>
      booth_integration_output_9_6, S0=>nx14668);
   ix3482 : mux21_ni port map ( Y=>nx3481, A0=>booth_integration_output_9_6, 
      A1=>nx762, S0=>nx14394);
   ix763 : mux21_ni port map ( Y=>nx762, A0=>neuron(6), A1=>
      booth_integration_output_9_7, S0=>nx14668);
   ix3472 : mux21_ni port map ( Y=>nx3471, A0=>booth_integration_output_9_7, 
      A1=>nx750, S0=>nx14658);
   ix751 : mux21_ni port map ( Y=>nx750, A0=>neuron(7), A1=>
      booth_integration_output_9_8, S0=>nx14668);
   ix3462 : mux21_ni port map ( Y=>nx3461, A0=>booth_integration_output_9_8, 
      A1=>nx738, S0=>nx14658);
   ix739 : mux21_ni port map ( Y=>nx738, A0=>neuron(8), A1=>
      booth_integration_output_9_9, S0=>nx14668);
   ix3452 : mux21_ni port map ( Y=>nx3451, A0=>booth_integration_output_9_9, 
      A1=>nx726, S0=>nx14658);
   ix727 : mux21_ni port map ( Y=>nx726, A0=>neuron(9), A1=>
      booth_integration_output_9_10, S0=>nx14668);
   ix3442 : mux21_ni port map ( Y=>nx3441, A0=>booth_integration_output_9_10, 
      A1=>nx714, S0=>nx14660);
   ix715 : mux21_ni port map ( Y=>nx714, A0=>neuron(10), A1=>
      booth_integration_output_9_11, S0=>nx14668);
   ix3432 : mux21_ni port map ( Y=>nx3431, A0=>booth_integration_output_9_11, 
      A1=>nx702, S0=>nx14660);
   ix703 : mux21_ni port map ( Y=>nx702, A0=>neuron(11), A1=>
      booth_integration_output_9_12, S0=>nx14668);
   ix3422 : mux21_ni port map ( Y=>nx3421, A0=>booth_integration_output_9_12, 
      A1=>nx690, S0=>nx14660);
   ix691 : mux21_ni port map ( Y=>nx690, A0=>neuron(12), A1=>
      booth_integration_output_9_13, S0=>nx14670);
   ix3412 : mux21_ni port map ( Y=>nx3411, A0=>booth_integration_output_9_13, 
      A1=>nx678, S0=>nx14660);
   ix679 : mux21_ni port map ( Y=>nx678, A0=>neuron(13), A1=>
      booth_integration_output_9_14, S0=>nx14670);
   ix3402 : mux21_ni port map ( Y=>nx3401, A0=>booth_integration_output_9_14, 
      A1=>nx666, S0=>nx14660);
   ix667 : mux21_ni port map ( Y=>nx666, A0=>neuron(14), A1=>
      booth_integration_output_9_15, S0=>nx14670);
   ix3392 : mux21 port map ( Y=>nx3391, A0=>nx9139, A1=>nx8668, S0=>nx14660
   );
   ix3042 : mux21_ni port map ( Y=>nx3041, A0=>
      booth_integrtaion_9_shift_Reg_count_0, A1=>nx14174, S0=>nx14612);
   ix3028 : and02 port map ( Y=>nx3027, A0=>nx14822, A1=>
      booth_integrtaion_9_shift_Reg_count_0);
   ix3222 : mux21_ni port map ( Y=>nx3221, A0=>
      booth_integrtaion_9_shift_Reg_count_9, A1=>nx14122, S0=>nx14612);
   ix3212 : mux21_ni port map ( Y=>nx3211, A0=>
      booth_integrtaion_9_shift_Reg_count_9, A1=>
      booth_integrtaion_9_shift_Reg_output_8, S0=>nx14660);
   ix3202 : mux21_ni port map ( Y=>nx3201, A0=>
      booth_integrtaion_9_shift_Reg_count_8, A1=>
      booth_integrtaion_9_shift_Reg_output_8, S0=>nx14612);
   ix3192 : mux21_ni port map ( Y=>nx3191, A0=>
      booth_integrtaion_9_shift_Reg_count_8, A1=>
      booth_integrtaion_9_shift_Reg_output_7, S0=>nx14662);
   ix3182 : mux21_ni port map ( Y=>nx3181, A0=>
      booth_integrtaion_9_shift_Reg_count_7, A1=>
      booth_integrtaion_9_shift_Reg_output_7, S0=>nx14612);
   ix3172 : mux21_ni port map ( Y=>nx3171, A0=>
      booth_integrtaion_9_shift_Reg_count_7, A1=>
      booth_integrtaion_9_shift_Reg_output_6, S0=>nx14662);
   ix3162 : mux21_ni port map ( Y=>nx3161, A0=>
      booth_integrtaion_9_shift_Reg_count_6, A1=>
      booth_integrtaion_9_shift_Reg_output_6, S0=>nx14612);
   ix3152 : mux21_ni port map ( Y=>nx3151, A0=>
      booth_integrtaion_9_shift_Reg_count_6, A1=>
      booth_integrtaion_9_shift_Reg_output_5, S0=>nx14662);
   ix3142 : mux21_ni port map ( Y=>nx3141, A0=>
      booth_integrtaion_9_shift_Reg_count_5, A1=>
      booth_integrtaion_9_shift_Reg_output_5, S0=>nx14612);
   ix3132 : mux21_ni port map ( Y=>nx3131, A0=>
      booth_integrtaion_9_shift_Reg_count_5, A1=>
      booth_integrtaion_9_shift_Reg_output_4, S0=>nx14662);
   ix3122 : mux21_ni port map ( Y=>nx3121, A0=>
      booth_integrtaion_9_shift_Reg_count_4, A1=>
      booth_integrtaion_9_shift_Reg_output_4, S0=>nx14614);
   ix3112 : mux21_ni port map ( Y=>nx3111, A0=>
      booth_integrtaion_9_shift_Reg_count_4, A1=>
      booth_integrtaion_9_shift_Reg_output_3, S0=>nx14662);
   ix3102 : mux21_ni port map ( Y=>nx3101, A0=>
      booth_integrtaion_9_shift_Reg_count_3, A1=>
      booth_integrtaion_9_shift_Reg_output_3, S0=>nx14614);
   ix3092 : mux21_ni port map ( Y=>nx3091, A0=>
      booth_integrtaion_9_shift_Reg_count_3, A1=>
      booth_integrtaion_9_shift_Reg_output_2, S0=>nx14662);
   ix3082 : mux21_ni port map ( Y=>nx3081, A0=>
      booth_integrtaion_9_shift_Reg_count_2, A1=>
      booth_integrtaion_9_shift_Reg_output_2, S0=>nx14614);
   ix3072 : mux21_ni port map ( Y=>nx3071, A0=>
      booth_integrtaion_9_shift_Reg_count_2, A1=>
      booth_integrtaion_9_shift_Reg_output_1, S0=>nx14662);
   ix3062 : mux21_ni port map ( Y=>nx3061, A0=>
      booth_integrtaion_9_shift_Reg_count_1, A1=>
      booth_integrtaion_9_shift_Reg_output_1, S0=>nx14614);
   ix3052 : mux21_ni port map ( Y=>nx3051, A0=>
      booth_integrtaion_9_shift_Reg_count_1, A1=>nx14174, S0=>nx14664);
   ix107 : and02 port map ( Y=>nx106, A0=>nx8777, A1=>
      booth_integration_output_9_0);
   ix8780 : or03 port map ( Y=>nx8779, A0=>nx8605, A1=>
      booth_integrtaion_9_shift_reg_output_0, A2=>nx14822);
   ix3382 : mux21_ni port map ( Y=>nx3381, A0=>
      booth_integrtaion_9_booth_output_16, A1=>nx636, S0=>nx14664);
   ix637 : nor02ii port map ( Y=>nx636, A0=>nx8791, A1=>nx14670);
   ix113 : nor02ii port map ( Y=>nx112, A0=>nx8769, A1=>
      booth_integrtaion_9_booth_output_16);
   ix631 : xor2 port map ( Y=>nx2805, A0=>nx8801, A1=>nx9133);
   ix619 : xor2 port map ( Y=>nx2807, A0=>nx8821, A1=>nx14400);
   ix3352 : mux21_ni port map ( Y=>nx3351, A0=>
      booth_integrtaion_9_booth_output_19, A1=>nx600, S0=>nx14664);
   ix601 : nor02ii port map ( Y=>nx600, A0=>nx8845, A1=>nx14670);
   ix8862 : nor02_2x port map ( Y=>nx102, A0=>nx8777, A1=>
      booth_integration_output_9_0);
   ix8866 : xor2 port map ( Y=>nx8865, A0=>nx8871, A1=>nx208);
   ix3332 : mux21_ni port map ( Y=>nx3331, A0=>
      booth_integrtaion_9_booth_output_21, A1=>nx576, S0=>nx14664);
   ix577 : nor02ii port map ( Y=>nx576, A0=>nx8893, A1=>nx14670);
   ix8906 : xor2 port map ( Y=>nx8905, A0=>nx8909, A1=>nx256);
   ix3312 : mux21_ni port map ( Y=>nx3311, A0=>
      booth_integrtaion_9_booth_output_23, A1=>nx552, S0=>nx14664);
   ix553 : nor02ii port map ( Y=>nx552, A0=>nx8929, A1=>nx14670);
   ix8942 : xor2 port map ( Y=>nx8941, A0=>nx8945, A1=>nx304);
   ix3292 : mux21_ni port map ( Y=>nx3291, A0=>
      booth_integrtaion_9_booth_output_25, A1=>nx528, S0=>nx14664);
   ix529 : nor02ii port map ( Y=>nx528, A0=>nx8965, A1=>nx14672);
   ix8980 : xor2 port map ( Y=>nx8979, A0=>nx8985, A1=>nx352);
   ix3272 : mux21_ni port map ( Y=>nx3271, A0=>
      booth_integrtaion_9_booth_output_27, A1=>nx504, S0=>nx14664);
   ix505 : nor02ii port map ( Y=>nx504, A0=>nx9011, A1=>nx14672);
   ix9028 : xor2 port map ( Y=>nx9027, A0=>nx9033, A1=>nx400);
   ix3252 : mux21_ni port map ( Y=>nx3251, A0=>
      booth_integrtaion_9_booth_output_29, A1=>nx480, S0=>nx14392);
   ix481 : nor02ii port map ( Y=>nx480, A0=>nx9059, A1=>nx14672);
   ix9076 : xor2 port map ( Y=>nx9075, A0=>nx9087, A1=>nx448);
   ix3242 : mux21_ni port map ( Y=>nx3241, A0=>
      booth_integrtaion_9_booth_output_31, A1=>nx468, S0=>nx14392);
   ix469 : nor02ii port map ( Y=>nx468, A0=>nx9083, A1=>nx14672);
   ix463 : xor2 port map ( Y=>nx462, A0=>nx9087, A1=>nx9101);
   ix649 : nor02ii port map ( Y=>nx648, A0=>nx112, A1=>nx14672);
   ix9176 : xor2 port map ( Y=>nx9175, A0=>nx9161, A1=>adderInput_9(2));
   ix9192 : xor2 port map ( Y=>nx9191, A0=>nx9157, A1=>adderInput_9(4));
   ix9208 : xor2 port map ( Y=>nx9207, A0=>nx9153, A1=>adderInput_9(6));
   ix9224 : xor2 port map ( Y=>nx9223, A0=>nx9149, A1=>adderInput_9(8));
   ix9240 : xor2 port map ( Y=>nx9239, A0=>nx9146, A1=>adderInput_9(10));
   ix9256 : xor2 port map ( Y=>nx9255, A0=>nx9143, A1=>adderInput_9(12));
   ix9272 : xor2 port map ( Y=>nx9271, A0=>nx9141, A1=>adderInput_9(14));
   ix9280 : xor2 port map ( Y=>nx9279, A0=>nx9139, A1=>adderInput_9(15));
   ix1977 : xor2 port map ( Y=>label_8(0), A0=>adderInput_8(0), A1=>
      booth_integration_output_8_0);
   ix4072 : mux21_ni port map ( Y=>nx4071, A0=>booth_integration_output_8_0, 
      A1=>nx1820, S0=>nx14416);
   ix1821 : mux21_ni port map ( Y=>nx1820, A0=>neuron(0), A1=>
      booth_integration_output_8_1, S0=>nx14682);
   ix4062 : mux21_ni port map ( Y=>nx4061, A0=>booth_integration_output_8_1, 
      A1=>nx1808, S0=>nx14416);
   ix1809 : mux21_ni port map ( Y=>nx1808, A0=>neuron(1), A1=>
      booth_integration_output_8_2, S0=>nx14682);
   ix4052 : mux21_ni port map ( Y=>nx4051, A0=>booth_integration_output_8_2, 
      A1=>nx1796, S0=>nx14416);
   ix1797 : mux21_ni port map ( Y=>nx1796, A0=>neuron(2), A1=>
      booth_integration_output_8_3, S0=>nx14682);
   ix4042 : mux21_ni port map ( Y=>nx4041, A0=>booth_integration_output_8_3, 
      A1=>nx1784, S0=>nx14416);
   ix1785 : mux21_ni port map ( Y=>nx1784, A0=>neuron(3), A1=>
      booth_integration_output_8_4, S0=>nx14682);
   ix4032 : mux21_ni port map ( Y=>nx4031, A0=>booth_integration_output_8_4, 
      A1=>nx1772, S0=>nx14416);
   ix1773 : mux21_ni port map ( Y=>nx1772, A0=>neuron(4), A1=>
      booth_integration_output_8_5, S0=>nx14682);
   ix4022 : mux21_ni port map ( Y=>nx4021, A0=>booth_integration_output_8_5, 
      A1=>nx1760, S0=>nx14416);
   ix1761 : mux21_ni port map ( Y=>nx1760, A0=>neuron(5), A1=>
      booth_integration_output_8_6, S0=>nx14684);
   ix4012 : mux21_ni port map ( Y=>nx4011, A0=>booth_integration_output_8_6, 
      A1=>nx1748, S0=>nx14416);
   ix1749 : mux21_ni port map ( Y=>nx1748, A0=>neuron(6), A1=>
      booth_integration_output_8_7, S0=>nx14684);
   ix4002 : mux21_ni port map ( Y=>nx4001, A0=>booth_integration_output_8_7, 
      A1=>nx1736, S0=>nx14674);
   ix1737 : mux21_ni port map ( Y=>nx1736, A0=>neuron(7), A1=>
      booth_integration_output_8_8, S0=>nx14684);
   ix3992 : mux21_ni port map ( Y=>nx3991, A0=>booth_integration_output_8_8, 
      A1=>nx1724, S0=>nx14674);
   ix1725 : mux21_ni port map ( Y=>nx1724, A0=>neuron(8), A1=>
      booth_integration_output_8_9, S0=>nx14684);
   ix3982 : mux21_ni port map ( Y=>nx3981, A0=>booth_integration_output_8_9, 
      A1=>nx1712, S0=>nx14674);
   ix1713 : mux21_ni port map ( Y=>nx1712, A0=>neuron(9), A1=>
      booth_integration_output_8_10, S0=>nx14684);
   ix3972 : mux21_ni port map ( Y=>nx3971, A0=>booth_integration_output_8_10, 
      A1=>nx1700, S0=>nx14676);
   ix1701 : mux21_ni port map ( Y=>nx1700, A0=>neuron(10), A1=>
      booth_integration_output_8_11, S0=>nx14684);
   ix3962 : mux21_ni port map ( Y=>nx3961, A0=>booth_integration_output_8_11, 
      A1=>nx1688, S0=>nx14676);
   ix1689 : mux21_ni port map ( Y=>nx1688, A0=>neuron(11), A1=>
      booth_integration_output_8_12, S0=>nx14684);
   ix3952 : mux21_ni port map ( Y=>nx3951, A0=>booth_integration_output_8_12, 
      A1=>nx1676, S0=>nx14676);
   ix1677 : mux21_ni port map ( Y=>nx1676, A0=>neuron(12), A1=>
      booth_integration_output_8_13, S0=>nx14686);
   ix3942 : mux21_ni port map ( Y=>nx3941, A0=>booth_integration_output_8_13, 
      A1=>nx1664, S0=>nx14676);
   ix1665 : mux21_ni port map ( Y=>nx1664, A0=>neuron(13), A1=>
      booth_integration_output_8_14, S0=>nx14686);
   ix3932 : mux21_ni port map ( Y=>nx3931, A0=>booth_integration_output_8_14, 
      A1=>nx1652, S0=>nx14676);
   ix1653 : mux21_ni port map ( Y=>nx1652, A0=>neuron(14), A1=>
      booth_integration_output_8_15, S0=>nx14686);
   ix3922 : mux21 port map ( Y=>nx3921, A0=>nx9811, A1=>nx9361, S0=>nx14676
   );
   ix3572 : mux21_ni port map ( Y=>nx3571, A0=>
      booth_integrtaion_8_shift_Reg_count_0, A1=>nx14196, S0=>nx14616);
   ix3558 : and02 port map ( Y=>nx3557, A0=>nx14826, A1=>
      booth_integrtaion_8_shift_Reg_count_0);
   ix3752 : mux21_ni port map ( Y=>nx3751, A0=>
      booth_integrtaion_8_shift_Reg_count_9, A1=>nx14182, S0=>nx14616);
   ix3742 : mux21_ni port map ( Y=>nx3741, A0=>
      booth_integrtaion_8_shift_Reg_count_9, A1=>
      booth_integrtaion_8_shift_Reg_output_8, S0=>nx14676);
   ix3732 : mux21_ni port map ( Y=>nx3731, A0=>
      booth_integrtaion_8_shift_Reg_count_8, A1=>
      booth_integrtaion_8_shift_Reg_output_8, S0=>nx14616);
   ix3722 : mux21_ni port map ( Y=>nx3721, A0=>
      booth_integrtaion_8_shift_Reg_count_8, A1=>
      booth_integrtaion_8_shift_Reg_output_7, S0=>nx14678);
   ix3712 : mux21_ni port map ( Y=>nx3711, A0=>
      booth_integrtaion_8_shift_Reg_count_7, A1=>
      booth_integrtaion_8_shift_Reg_output_7, S0=>nx14616);
   ix3702 : mux21_ni port map ( Y=>nx3701, A0=>
      booth_integrtaion_8_shift_Reg_count_7, A1=>
      booth_integrtaion_8_shift_Reg_output_6, S0=>nx14678);
   ix3692 : mux21_ni port map ( Y=>nx3691, A0=>
      booth_integrtaion_8_shift_Reg_count_6, A1=>
      booth_integrtaion_8_shift_Reg_output_6, S0=>nx14616);
   ix3682 : mux21_ni port map ( Y=>nx3681, A0=>
      booth_integrtaion_8_shift_Reg_count_6, A1=>
      booth_integrtaion_8_shift_Reg_output_5, S0=>nx14678);
   ix3672 : mux21_ni port map ( Y=>nx3671, A0=>
      booth_integrtaion_8_shift_Reg_count_5, A1=>
      booth_integrtaion_8_shift_Reg_output_5, S0=>nx14616);
   ix3662 : mux21_ni port map ( Y=>nx3661, A0=>
      booth_integrtaion_8_shift_Reg_count_5, A1=>
      booth_integrtaion_8_shift_Reg_output_4, S0=>nx14678);
   ix3652 : mux21_ni port map ( Y=>nx3651, A0=>
      booth_integrtaion_8_shift_Reg_count_4, A1=>
      booth_integrtaion_8_shift_Reg_output_4, S0=>nx14618);
   ix3642 : mux21_ni port map ( Y=>nx3641, A0=>
      booth_integrtaion_8_shift_Reg_count_4, A1=>
      booth_integrtaion_8_shift_Reg_output_3, S0=>nx14678);
   ix3632 : mux21_ni port map ( Y=>nx3631, A0=>
      booth_integrtaion_8_shift_Reg_count_3, A1=>
      booth_integrtaion_8_shift_Reg_output_3, S0=>nx14618);
   ix3622 : mux21_ni port map ( Y=>nx3621, A0=>
      booth_integrtaion_8_shift_Reg_count_3, A1=>
      booth_integrtaion_8_shift_Reg_output_2, S0=>nx14678);
   ix3612 : mux21_ni port map ( Y=>nx3611, A0=>
      booth_integrtaion_8_shift_Reg_count_2, A1=>
      booth_integrtaion_8_shift_Reg_output_2, S0=>nx14618);
   ix3602 : mux21_ni port map ( Y=>nx3601, A0=>
      booth_integrtaion_8_shift_Reg_count_2, A1=>
      booth_integrtaion_8_shift_Reg_output_1, S0=>nx14678);
   ix3592 : mux21_ni port map ( Y=>nx3591, A0=>
      booth_integrtaion_8_shift_Reg_count_1, A1=>
      booth_integrtaion_8_shift_Reg_output_1, S0=>nx14618);
   ix3582 : mux21_ni port map ( Y=>nx3581, A0=>
      booth_integrtaion_8_shift_Reg_count_1, A1=>nx14196, S0=>nx14680);
   ix1093 : and02 port map ( Y=>nx1092, A0=>nx9453, A1=>
      booth_integration_output_8_0);
   ix9456 : or03 port map ( Y=>nx9455, A0=>nx9283, A1=>
      booth_integrtaion_8_shift_reg_output_0, A2=>nx14826);
   ix3912 : mux21_ni port map ( Y=>nx3911, A0=>
      booth_integrtaion_8_booth_output_16, A1=>nx1622, S0=>nx14680);
   ix1623 : nor02ii port map ( Y=>nx1622, A0=>nx9466, A1=>nx14686);
   ix1099 : nor02ii port map ( Y=>nx1098, A0=>nx9447, A1=>
      booth_integrtaion_8_booth_output_16);
   ix1617 : xor2 port map ( Y=>nx2831, A0=>nx9475, A1=>nx9805);
   ix1605 : xor2 port map ( Y=>nx2833, A0=>nx9492, A1=>nx14422);
   ix3882 : mux21_ni port map ( Y=>nx3881, A0=>
      booth_integrtaion_8_booth_output_19, A1=>nx1586, S0=>nx14680);
   ix1587 : nor02ii port map ( Y=>nx1586, A0=>nx9513, A1=>nx14686);
   ix9530 : nor02_2x port map ( Y=>nx1088, A0=>nx9453, A1=>
      booth_integration_output_8_0);
   ix9533 : xor2 port map ( Y=>nx9532, A0=>nx9537, A1=>nx1194);
   ix3862 : mux21_ni port map ( Y=>nx3861, A0=>
      booth_integrtaion_8_booth_output_21, A1=>nx1562, S0=>nx14680);
   ix1563 : nor02ii port map ( Y=>nx1562, A0=>nx9558, A1=>nx14686);
   ix9574 : xor2 port map ( Y=>nx9573, A0=>nx9579, A1=>nx1242);
   ix3842 : mux21_ni port map ( Y=>nx3841, A0=>
      booth_integrtaion_8_booth_output_23, A1=>nx1538, S0=>nx14680);
   ix1539 : nor02ii port map ( Y=>nx1538, A0=>nx9603, A1=>nx14686);
   ix9619 : xor2 port map ( Y=>nx9618, A0=>nx9623, A1=>nx1290);
   ix3822 : mux21_ni port map ( Y=>nx3821, A0=>
      booth_integrtaion_8_booth_output_25, A1=>nx1514, S0=>nx14680);
   ix1515 : nor02ii port map ( Y=>nx1514, A0=>nx9645, A1=>nx14688);
   ix9660 : xor2 port map ( Y=>nx9659, A0=>nx9664, A1=>nx1338);
   ix3802 : mux21_ni port map ( Y=>nx3801, A0=>
      booth_integrtaion_8_booth_output_27, A1=>nx1490, S0=>nx14680);
   ix1491 : nor02ii port map ( Y=>nx1490, A0=>nx9688, A1=>nx14688);
   ix9703 : xor2 port map ( Y=>nx9702, A0=>nx9707, A1=>nx1386);
   ix3782 : mux21_ni port map ( Y=>nx3781, A0=>
      booth_integrtaion_8_booth_output_29, A1=>nx1466, S0=>nx14414);
   ix1467 : nor02ii port map ( Y=>nx1466, A0=>nx9731, A1=>nx14688);
   ix9748 : xor2 port map ( Y=>nx9747, A0=>nx9759, A1=>nx1434);
   ix3772 : mux21_ni port map ( Y=>nx3771, A0=>
      booth_integrtaion_8_booth_output_31, A1=>nx1454, S0=>nx14414);
   ix1455 : nor02ii port map ( Y=>nx1454, A0=>nx9755, A1=>nx14688);
   ix1449 : xor2 port map ( Y=>nx1448, A0=>nx9759, A1=>nx9773);
   ix1635 : nor02ii port map ( Y=>nx1634, A0=>nx1098, A1=>nx14688);
   ix9848 : xor2 port map ( Y=>nx9847, A0=>nx9833, A1=>adderInput_8(2));
   ix9864 : xor2 port map ( Y=>nx9863, A0=>nx9831, A1=>adderInput_8(4));
   ix9878 : xor2 port map ( Y=>nx9877, A0=>nx9829, A1=>adderInput_8(6));
   ix9890 : xor2 port map ( Y=>nx9889, A0=>nx9825, A1=>adderInput_8(8));
   ix9902 : xor2 port map ( Y=>nx9901, A0=>nx9821, A1=>adderInput_8(10));
   ix9914 : xor2 port map ( Y=>nx9913, A0=>nx9817, A1=>adderInput_8(12));
   ix9926 : xor2 port map ( Y=>nx9925, A0=>nx9813, A1=>adderInput_8(14));
   ix9932 : xor2 port map ( Y=>nx9931, A0=>nx9811, A1=>adderInput_8(15));
   ix2963 : xor2 port map ( Y=>label_7(0), A0=>adderInput_7(0), A1=>
      booth_integration_output_7_0);
   ix4602 : mux21_ni port map ( Y=>nx4601, A0=>booth_integration_output_7_0, 
      A1=>nx2806, S0=>nx14438);
   ix2807 : mux21_ni port map ( Y=>nx2806, A0=>neuron(0), A1=>
      booth_integration_output_7_1, S0=>nx14698);
   ix4592 : mux21_ni port map ( Y=>nx4591, A0=>booth_integration_output_7_1, 
      A1=>nx2794, S0=>nx14438);
   ix2795 : mux21_ni port map ( Y=>nx2794, A0=>neuron(1), A1=>
      booth_integration_output_7_2, S0=>nx14698);
   ix4582 : mux21_ni port map ( Y=>nx4581, A0=>booth_integration_output_7_2, 
      A1=>nx2782, S0=>nx14438);
   ix2783 : mux21_ni port map ( Y=>nx2782, A0=>neuron(2), A1=>
      booth_integration_output_7_3, S0=>nx14698);
   ix4572 : mux21_ni port map ( Y=>nx4571, A0=>booth_integration_output_7_3, 
      A1=>nx2770, S0=>nx14438);
   ix2771 : mux21_ni port map ( Y=>nx2770, A0=>neuron(3), A1=>
      booth_integration_output_7_4, S0=>nx14698);
   ix4562 : mux21_ni port map ( Y=>nx4561, A0=>booth_integration_output_7_4, 
      A1=>nx2758, S0=>nx14438);
   ix2759 : mux21_ni port map ( Y=>nx2758, A0=>neuron(4), A1=>
      booth_integration_output_7_5, S0=>nx14698);
   ix4552 : mux21_ni port map ( Y=>nx4551, A0=>booth_integration_output_7_5, 
      A1=>nx2746, S0=>nx14438);
   ix2747 : mux21_ni port map ( Y=>nx2746, A0=>neuron(5), A1=>
      booth_integration_output_7_6, S0=>nx14700);
   ix4542 : mux21_ni port map ( Y=>nx4541, A0=>booth_integration_output_7_6, 
      A1=>nx2734, S0=>nx14438);
   ix2735 : mux21_ni port map ( Y=>nx2734, A0=>neuron(6), A1=>
      booth_integration_output_7_7, S0=>nx14700);
   ix4532 : mux21_ni port map ( Y=>nx4531, A0=>booth_integration_output_7_7, 
      A1=>nx2722, S0=>nx14690);
   ix2723 : mux21_ni port map ( Y=>nx2722, A0=>neuron(7), A1=>
      booth_integration_output_7_8, S0=>nx14700);
   ix4522 : mux21_ni port map ( Y=>nx4521, A0=>booth_integration_output_7_8, 
      A1=>nx2710, S0=>nx14690);
   ix2711 : mux21_ni port map ( Y=>nx2710, A0=>neuron(8), A1=>
      booth_integration_output_7_9, S0=>nx14700);
   ix4512 : mux21_ni port map ( Y=>nx4511, A0=>booth_integration_output_7_9, 
      A1=>nx2698, S0=>nx14690);
   ix2699 : mux21_ni port map ( Y=>nx2698, A0=>neuron(9), A1=>
      booth_integration_output_7_10, S0=>nx14700);
   ix4502 : mux21_ni port map ( Y=>nx4501, A0=>booth_integration_output_7_10, 
      A1=>nx2686, S0=>nx14692);
   ix2687 : mux21_ni port map ( Y=>nx2686, A0=>neuron(10), A1=>
      booth_integration_output_7_11, S0=>nx14700);
   ix4492 : mux21_ni port map ( Y=>nx4491, A0=>booth_integration_output_7_11, 
      A1=>nx2674, S0=>nx14692);
   ix2675 : mux21_ni port map ( Y=>nx2674, A0=>neuron(11), A1=>
      booth_integration_output_7_12, S0=>nx14700);
   ix4482 : mux21_ni port map ( Y=>nx4481, A0=>booth_integration_output_7_12, 
      A1=>nx2662, S0=>nx14692);
   ix2663 : mux21_ni port map ( Y=>nx2662, A0=>neuron(12), A1=>
      booth_integration_output_7_13, S0=>nx14702);
   ix4472 : mux21_ni port map ( Y=>nx4471, A0=>booth_integration_output_7_13, 
      A1=>nx2650, S0=>nx14692);
   ix2651 : mux21_ni port map ( Y=>nx2650, A0=>neuron(13), A1=>
      booth_integration_output_7_14, S0=>nx14702);
   ix4462 : mux21_ni port map ( Y=>nx4461, A0=>booth_integration_output_7_14, 
      A1=>nx2638, S0=>nx14692);
   ix2639 : mux21_ni port map ( Y=>nx2638, A0=>neuron(14), A1=>
      booth_integration_output_7_15, S0=>nx14702);
   ix4452 : mux21 port map ( Y=>nx4451, A0=>nx10351, A1=>nx9982, S0=>nx14692
   );
   ix4102 : mux21_ni port map ( Y=>nx4101, A0=>
      booth_integrtaion_7_shift_Reg_count_0, A1=>nx14218, S0=>nx14620);
   ix4088 : and02 port map ( Y=>nx4087, A0=>nx14830, A1=>
      booth_integrtaion_7_shift_Reg_count_0);
   ix4282 : mux21_ni port map ( Y=>nx4281, A0=>
      booth_integrtaion_7_shift_Reg_count_9, A1=>nx14204, S0=>nx14620);
   ix4272 : mux21_ni port map ( Y=>nx4271, A0=>
      booth_integrtaion_7_shift_Reg_count_9, A1=>
      booth_integrtaion_7_shift_Reg_output_8, S0=>nx14692);
   ix4262 : mux21_ni port map ( Y=>nx4261, A0=>
      booth_integrtaion_7_shift_Reg_count_8, A1=>
      booth_integrtaion_7_shift_Reg_output_8, S0=>nx14620);
   ix4252 : mux21_ni port map ( Y=>nx4251, A0=>
      booth_integrtaion_7_shift_Reg_count_8, A1=>
      booth_integrtaion_7_shift_Reg_output_7, S0=>nx14694);
   ix4242 : mux21_ni port map ( Y=>nx4241, A0=>
      booth_integrtaion_7_shift_Reg_count_7, A1=>
      booth_integrtaion_7_shift_Reg_output_7, S0=>nx14620);
   ix4232 : mux21_ni port map ( Y=>nx4231, A0=>
      booth_integrtaion_7_shift_Reg_count_7, A1=>
      booth_integrtaion_7_shift_Reg_output_6, S0=>nx14694);
   ix4222 : mux21_ni port map ( Y=>nx4221, A0=>
      booth_integrtaion_7_shift_Reg_count_6, A1=>
      booth_integrtaion_7_shift_Reg_output_6, S0=>nx14620);
   ix4212 : mux21_ni port map ( Y=>nx4211, A0=>
      booth_integrtaion_7_shift_Reg_count_6, A1=>
      booth_integrtaion_7_shift_Reg_output_5, S0=>nx14694);
   ix4202 : mux21_ni port map ( Y=>nx4201, A0=>
      booth_integrtaion_7_shift_Reg_count_5, A1=>
      booth_integrtaion_7_shift_Reg_output_5, S0=>nx14620);
   ix4192 : mux21_ni port map ( Y=>nx4191, A0=>
      booth_integrtaion_7_shift_Reg_count_5, A1=>
      booth_integrtaion_7_shift_Reg_output_4, S0=>nx14694);
   ix4182 : mux21_ni port map ( Y=>nx4181, A0=>
      booth_integrtaion_7_shift_Reg_count_4, A1=>
      booth_integrtaion_7_shift_Reg_output_4, S0=>nx14622);
   ix4172 : mux21_ni port map ( Y=>nx4171, A0=>
      booth_integrtaion_7_shift_Reg_count_4, A1=>
      booth_integrtaion_7_shift_Reg_output_3, S0=>nx14694);
   ix4162 : mux21_ni port map ( Y=>nx4161, A0=>
      booth_integrtaion_7_shift_Reg_count_3, A1=>
      booth_integrtaion_7_shift_Reg_output_3, S0=>nx14622);
   ix4152 : mux21_ni port map ( Y=>nx4151, A0=>
      booth_integrtaion_7_shift_Reg_count_3, A1=>
      booth_integrtaion_7_shift_Reg_output_2, S0=>nx14694);
   ix4142 : mux21_ni port map ( Y=>nx4141, A0=>
      booth_integrtaion_7_shift_Reg_count_2, A1=>
      booth_integrtaion_7_shift_Reg_output_2, S0=>nx14622);
   ix4132 : mux21_ni port map ( Y=>nx4131, A0=>
      booth_integrtaion_7_shift_Reg_count_2, A1=>
      booth_integrtaion_7_shift_Reg_output_1, S0=>nx14694);
   ix4122 : mux21_ni port map ( Y=>nx4121, A0=>
      booth_integrtaion_7_shift_Reg_count_1, A1=>
      booth_integrtaion_7_shift_Reg_output_1, S0=>nx14622);
   ix4112 : mux21_ni port map ( Y=>nx4111, A0=>
      booth_integrtaion_7_shift_Reg_count_1, A1=>nx14218, S0=>nx14696);
   ix2079 : and02 port map ( Y=>nx2078, A0=>nx10055, A1=>
      booth_integration_output_7_0);
   ix10058 : or03 port map ( Y=>nx10057, A0=>nx9934, A1=>
      booth_integrtaion_7_shift_reg_output_0, A2=>nx14830);
   ix4442 : mux21_ni port map ( Y=>nx4441, A0=>
      booth_integrtaion_7_booth_output_16, A1=>nx2608, S0=>nx14696);
   ix2609 : nor02ii port map ( Y=>nx2608, A0=>nx10065, A1=>nx14702);
   ix2085 : nor02ii port map ( Y=>nx2084, A0=>nx10050, A1=>
      booth_integrtaion_7_booth_output_16);
   ix2603 : xor2 port map ( Y=>nx2861, A0=>nx10071, A1=>nx10347);
   ix2591 : xor2 port map ( Y=>nx2863, A0=>nx10085, A1=>nx14444);
   ix4412 : mux21_ni port map ( Y=>nx4411, A0=>
      booth_integrtaion_7_booth_output_19, A1=>nx2572, S0=>nx14696);
   ix2573 : nor02ii port map ( Y=>nx2572, A0=>nx10103, A1=>nx14702);
   ix10117 : nor02_2x port map ( Y=>nx2074, A0=>nx10055, A1=>
      booth_integration_output_7_0);
   ix10120 : xor2 port map ( Y=>nx10119, A0=>nx10123, A1=>nx2180);
   ix4392 : mux21_ni port map ( Y=>nx4391, A0=>
      booth_integrtaion_7_booth_output_21, A1=>nx2548, S0=>nx14696);
   ix2549 : nor02ii port map ( Y=>nx2548, A0=>nx10143, A1=>nx14702);
   ix10156 : xor2 port map ( Y=>nx10155, A0=>nx10159, A1=>nx2228);
   ix4372 : mux21_ni port map ( Y=>nx4371, A0=>
      booth_integrtaion_7_booth_output_23, A1=>nx2524, S0=>nx14696);
   ix2525 : nor02ii port map ( Y=>nx2524, A0=>nx10179, A1=>nx14702);
   ix10192 : xor2 port map ( Y=>nx10191, A0=>nx10195, A1=>nx2276);
   ix4352 : mux21_ni port map ( Y=>nx4351, A0=>
      booth_integrtaion_7_booth_output_25, A1=>nx2500, S0=>nx14696);
   ix2501 : nor02ii port map ( Y=>nx2500, A0=>nx10215, A1=>nx14704);
   ix10228 : xor2 port map ( Y=>nx10227, A0=>nx10231, A1=>nx2324);
   ix4332 : mux21_ni port map ( Y=>nx4331, A0=>
      booth_integrtaion_7_booth_output_27, A1=>nx2476, S0=>nx14696);
   ix2477 : nor02ii port map ( Y=>nx2476, A0=>nx10251, A1=>nx14704);
   ix10264 : xor2 port map ( Y=>nx10263, A0=>nx10267, A1=>nx2372);
   ix4312 : mux21_ni port map ( Y=>nx4311, A0=>
      booth_integrtaion_7_booth_output_29, A1=>nx2452, S0=>nx14436);
   ix2453 : nor02ii port map ( Y=>nx2452, A0=>nx10287, A1=>nx14704);
   ix10300 : xor2 port map ( Y=>nx10299, A0=>nx10307, A1=>nx2420);
   ix4302 : mux21_ni port map ( Y=>nx4301, A0=>
      booth_integrtaion_7_booth_output_31, A1=>nx2440, S0=>nx14436);
   ix2441 : nor02ii port map ( Y=>nx2440, A0=>nx10304, A1=>nx14704);
   ix2435 : xor2 port map ( Y=>nx2434, A0=>nx10307, A1=>nx10319);
   ix2621 : nor02ii port map ( Y=>nx2620, A0=>nx2084, A1=>nx14704);
   ix10377 : xor2 port map ( Y=>nx10376, A0=>nx10365, A1=>adderInput_7(2));
   ix10389 : xor2 port map ( Y=>nx10388, A0=>nx10363, A1=>adderInput_7(4));
   ix10401 : xor2 port map ( Y=>nx10400, A0=>nx10361, A1=>adderInput_7(6));
   ix10413 : xor2 port map ( Y=>nx10412, A0=>nx10359, A1=>adderInput_7(8));
   ix10425 : xor2 port map ( Y=>nx10424, A0=>nx10357, A1=>adderInput_7(10));
   ix10437 : xor2 port map ( Y=>nx10436, A0=>nx10355, A1=>adderInput_7(12));
   ix10449 : xor2 port map ( Y=>nx10448, A0=>nx10353, A1=>adderInput_7(14));
   ix10455 : xor2 port map ( Y=>nx10454, A0=>nx10351, A1=>adderInput_7(15));
   ix3949 : xor2 port map ( Y=>label_6(0), A0=>adderInput_6(0), A1=>
      booth_integration_output_6_0);
   ix5132 : mux21_ni port map ( Y=>nx5131, A0=>booth_integration_output_6_0, 
      A1=>nx3792, S0=>nx14460);
   ix3793 : mux21_ni port map ( Y=>nx3792, A0=>neuron(0), A1=>
      booth_integration_output_6_1, S0=>nx14714);
   ix5122 : mux21_ni port map ( Y=>nx5121, A0=>booth_integration_output_6_1, 
      A1=>nx3780, S0=>nx14460);
   ix3781 : mux21_ni port map ( Y=>nx3780, A0=>neuron(1), A1=>
      booth_integration_output_6_2, S0=>nx14714);
   ix5112 : mux21_ni port map ( Y=>nx5111, A0=>booth_integration_output_6_2, 
      A1=>nx3768, S0=>nx14460);
   ix3769 : mux21_ni port map ( Y=>nx3768, A0=>neuron(2), A1=>
      booth_integration_output_6_3, S0=>nx14714);
   ix5102 : mux21_ni port map ( Y=>nx5101, A0=>booth_integration_output_6_3, 
      A1=>nx3756, S0=>nx14460);
   ix3757 : mux21_ni port map ( Y=>nx3756, A0=>neuron(3), A1=>
      booth_integration_output_6_4, S0=>nx14714);
   ix5092 : mux21_ni port map ( Y=>nx5091, A0=>booth_integration_output_6_4, 
      A1=>nx3744, S0=>nx14460);
   ix3745 : mux21_ni port map ( Y=>nx3744, A0=>neuron(4), A1=>
      booth_integration_output_6_5, S0=>nx14714);
   ix5082 : mux21_ni port map ( Y=>nx5081, A0=>booth_integration_output_6_5, 
      A1=>nx3732, S0=>nx14460);
   ix3733 : mux21_ni port map ( Y=>nx3732, A0=>neuron(5), A1=>
      booth_integration_output_6_6, S0=>nx14716);
   ix5072 : mux21_ni port map ( Y=>nx5071, A0=>booth_integration_output_6_6, 
      A1=>nx3720, S0=>nx14460);
   ix3721 : mux21_ni port map ( Y=>nx3720, A0=>neuron(6), A1=>
      booth_integration_output_6_7, S0=>nx14716);
   ix5062 : mux21_ni port map ( Y=>nx5061, A0=>booth_integration_output_6_7, 
      A1=>nx3708, S0=>nx14706);
   ix3709 : mux21_ni port map ( Y=>nx3708, A0=>neuron(7), A1=>
      booth_integration_output_6_8, S0=>nx14716);
   ix5052 : mux21_ni port map ( Y=>nx5051, A0=>booth_integration_output_6_8, 
      A1=>nx3696, S0=>nx14706);
   ix3697 : mux21_ni port map ( Y=>nx3696, A0=>neuron(8), A1=>
      booth_integration_output_6_9, S0=>nx14716);
   ix5042 : mux21_ni port map ( Y=>nx5041, A0=>booth_integration_output_6_9, 
      A1=>nx3684, S0=>nx14706);
   ix3685 : mux21_ni port map ( Y=>nx3684, A0=>neuron(9), A1=>
      booth_integration_output_6_10, S0=>nx14716);
   ix5032 : mux21_ni port map ( Y=>nx5031, A0=>booth_integration_output_6_10, 
      A1=>nx3672, S0=>nx14708);
   ix3673 : mux21_ni port map ( Y=>nx3672, A0=>neuron(10), A1=>
      booth_integration_output_6_11, S0=>nx14716);
   ix5022 : mux21_ni port map ( Y=>nx5021, A0=>booth_integration_output_6_11, 
      A1=>nx3660, S0=>nx14708);
   ix3661 : mux21_ni port map ( Y=>nx3660, A0=>neuron(11), A1=>
      booth_integration_output_6_12, S0=>nx14716);
   ix5012 : mux21_ni port map ( Y=>nx5011, A0=>booth_integration_output_6_12, 
      A1=>nx3648, S0=>nx14708);
   ix3649 : mux21_ni port map ( Y=>nx3648, A0=>neuron(12), A1=>
      booth_integration_output_6_13, S0=>nx14718);
   ix5002 : mux21_ni port map ( Y=>nx5001, A0=>booth_integration_output_6_13, 
      A1=>nx3636, S0=>nx14708);
   ix3637 : mux21_ni port map ( Y=>nx3636, A0=>neuron(13), A1=>
      booth_integration_output_6_14, S0=>nx14718);
   ix4992 : mux21_ni port map ( Y=>nx4991, A0=>booth_integration_output_6_14, 
      A1=>nx3624, S0=>nx14708);
   ix3625 : mux21_ni port map ( Y=>nx3624, A0=>neuron(14), A1=>
      booth_integration_output_6_15, S0=>nx14718);
   ix4982 : mux21 port map ( Y=>nx4981, A0=>nx10874, A1=>nx10505, S0=>
      nx14708);
   ix4632 : mux21_ni port map ( Y=>nx4631, A0=>
      booth_integrtaion_6_shift_Reg_count_0, A1=>nx14240, S0=>nx14624);
   ix4618 : and02 port map ( Y=>nx4617, A0=>nx14834, A1=>
      booth_integrtaion_6_shift_Reg_count_0);
   ix4812 : mux21_ni port map ( Y=>nx4811, A0=>
      booth_integrtaion_6_shift_Reg_count_9, A1=>nx14226, S0=>nx14624);
   ix4802 : mux21_ni port map ( Y=>nx4801, A0=>
      booth_integrtaion_6_shift_Reg_count_9, A1=>
      booth_integrtaion_6_shift_Reg_output_8, S0=>nx14708);
   ix4792 : mux21_ni port map ( Y=>nx4791, A0=>
      booth_integrtaion_6_shift_Reg_count_8, A1=>
      booth_integrtaion_6_shift_Reg_output_8, S0=>nx14624);
   ix4782 : mux21_ni port map ( Y=>nx4781, A0=>
      booth_integrtaion_6_shift_Reg_count_8, A1=>
      booth_integrtaion_6_shift_Reg_output_7, S0=>nx14710);
   ix4772 : mux21_ni port map ( Y=>nx4771, A0=>
      booth_integrtaion_6_shift_Reg_count_7, A1=>
      booth_integrtaion_6_shift_Reg_output_7, S0=>nx14624);
   ix4762 : mux21_ni port map ( Y=>nx4761, A0=>
      booth_integrtaion_6_shift_Reg_count_7, A1=>
      booth_integrtaion_6_shift_Reg_output_6, S0=>nx14710);
   ix4752 : mux21_ni port map ( Y=>nx4751, A0=>
      booth_integrtaion_6_shift_Reg_count_6, A1=>
      booth_integrtaion_6_shift_Reg_output_6, S0=>nx14624);
   ix4742 : mux21_ni port map ( Y=>nx4741, A0=>
      booth_integrtaion_6_shift_Reg_count_6, A1=>
      booth_integrtaion_6_shift_Reg_output_5, S0=>nx14710);
   ix4732 : mux21_ni port map ( Y=>nx4731, A0=>
      booth_integrtaion_6_shift_Reg_count_5, A1=>
      booth_integrtaion_6_shift_Reg_output_5, S0=>nx14624);
   ix4722 : mux21_ni port map ( Y=>nx4721, A0=>
      booth_integrtaion_6_shift_Reg_count_5, A1=>
      booth_integrtaion_6_shift_Reg_output_4, S0=>nx14710);
   ix4712 : mux21_ni port map ( Y=>nx4711, A0=>
      booth_integrtaion_6_shift_Reg_count_4, A1=>
      booth_integrtaion_6_shift_Reg_output_4, S0=>nx14626);
   ix4702 : mux21_ni port map ( Y=>nx4701, A0=>
      booth_integrtaion_6_shift_Reg_count_4, A1=>
      booth_integrtaion_6_shift_Reg_output_3, S0=>nx14710);
   ix4692 : mux21_ni port map ( Y=>nx4691, A0=>
      booth_integrtaion_6_shift_Reg_count_3, A1=>
      booth_integrtaion_6_shift_Reg_output_3, S0=>nx14626);
   ix4682 : mux21_ni port map ( Y=>nx4681, A0=>
      booth_integrtaion_6_shift_Reg_count_3, A1=>
      booth_integrtaion_6_shift_Reg_output_2, S0=>nx14710);
   ix4672 : mux21_ni port map ( Y=>nx4671, A0=>
      booth_integrtaion_6_shift_Reg_count_2, A1=>
      booth_integrtaion_6_shift_Reg_output_2, S0=>nx14626);
   ix4662 : mux21_ni port map ( Y=>nx4661, A0=>
      booth_integrtaion_6_shift_Reg_count_2, A1=>
      booth_integrtaion_6_shift_Reg_output_1, S0=>nx14710);
   ix4652 : mux21_ni port map ( Y=>nx4651, A0=>
      booth_integrtaion_6_shift_Reg_count_1, A1=>
      booth_integrtaion_6_shift_Reg_output_1, S0=>nx14626);
   ix4642 : mux21_ni port map ( Y=>nx4641, A0=>
      booth_integrtaion_6_shift_Reg_count_1, A1=>nx14240, S0=>nx14712);
   ix3065 : and02 port map ( Y=>nx3064, A0=>nx10578, A1=>
      booth_integration_output_6_0);
   ix10581 : or03 port map ( Y=>nx10580, A0=>nx10457, A1=>
      booth_integrtaion_6_shift_reg_output_0, A2=>nx14834);
   ix4972 : mux21_ni port map ( Y=>nx4971, A0=>
      booth_integrtaion_6_booth_output_16, A1=>nx3594, S0=>nx14712);
   ix3595 : nor02ii port map ( Y=>nx3594, A0=>nx10588, A1=>nx14718);
   ix3071 : nor02ii port map ( Y=>nx3070, A0=>nx10573, A1=>
      booth_integrtaion_6_booth_output_16);
   ix3589 : xor2 port map ( Y=>nx2891, A0=>nx10594, A1=>nx10870);
   ix3577 : xor2 port map ( Y=>nx2893, A0=>nx10608, A1=>nx14466);
   ix4942 : mux21_ni port map ( Y=>nx4941, A0=>
      booth_integrtaion_6_booth_output_19, A1=>nx3558, S0=>nx14712);
   ix3559 : nor02ii port map ( Y=>nx3558, A0=>nx10626, A1=>nx14718);
   ix10640 : nor02_2x port map ( Y=>nx3060, A0=>nx10578, A1=>
      booth_integration_output_6_0);
   ix10643 : xor2 port map ( Y=>nx10642, A0=>nx10646, A1=>nx3166);
   ix4922 : mux21_ni port map ( Y=>nx4921, A0=>
      booth_integrtaion_6_booth_output_21, A1=>nx3534, S0=>nx14712);
   ix3535 : nor02ii port map ( Y=>nx3534, A0=>nx10666, A1=>nx14718);
   ix10679 : xor2 port map ( Y=>nx10678, A0=>nx10682, A1=>nx3214);
   ix4902 : mux21_ni port map ( Y=>nx4901, A0=>
      booth_integrtaion_6_booth_output_23, A1=>nx3510, S0=>nx14712);
   ix3511 : nor02ii port map ( Y=>nx3510, A0=>nx10702, A1=>nx14718);
   ix10715 : xor2 port map ( Y=>nx10714, A0=>nx10718, A1=>nx3262);
   ix4882 : mux21_ni port map ( Y=>nx4881, A0=>
      booth_integrtaion_6_booth_output_25, A1=>nx3486, S0=>nx14712);
   ix3487 : nor02ii port map ( Y=>nx3486, A0=>nx10738, A1=>nx14720);
   ix10751 : xor2 port map ( Y=>nx10750, A0=>nx10754, A1=>nx3310);
   ix4862 : mux21_ni port map ( Y=>nx4861, A0=>
      booth_integrtaion_6_booth_output_27, A1=>nx3462, S0=>nx14712);
   ix3463 : nor02ii port map ( Y=>nx3462, A0=>nx10774, A1=>nx14720);
   ix10787 : xor2 port map ( Y=>nx10786, A0=>nx10790, A1=>nx3358);
   ix4842 : mux21_ni port map ( Y=>nx4841, A0=>
      booth_integrtaion_6_booth_output_29, A1=>nx3438, S0=>nx14458);
   ix3439 : nor02ii port map ( Y=>nx3438, A0=>nx10810, A1=>nx14720);
   ix10823 : xor2 port map ( Y=>nx10822, A0=>nx10830, A1=>nx3406);
   ix4832 : mux21_ni port map ( Y=>nx4831, A0=>
      booth_integrtaion_6_booth_output_31, A1=>nx3426, S0=>nx14458);
   ix3427 : nor02ii port map ( Y=>nx3426, A0=>nx10827, A1=>nx14720);
   ix3421 : xor2 port map ( Y=>nx3420, A0=>nx10830, A1=>nx10842);
   ix3607 : nor02ii port map ( Y=>nx3606, A0=>nx3070, A1=>nx14720);
   ix10900 : xor2 port map ( Y=>nx10899, A0=>nx10888, A1=>adderInput_6(2));
   ix10912 : xor2 port map ( Y=>nx10911, A0=>nx10886, A1=>adderInput_6(4));
   ix10924 : xor2 port map ( Y=>nx10923, A0=>nx10884, A1=>adderInput_6(6));
   ix10936 : xor2 port map ( Y=>nx10935, A0=>nx10882, A1=>adderInput_6(8));
   ix10948 : xor2 port map ( Y=>nx10947, A0=>nx10880, A1=>adderInput_6(10));
   ix10960 : xor2 port map ( Y=>nx10959, A0=>nx10878, A1=>adderInput_6(12));
   ix10972 : xor2 port map ( Y=>nx10971, A0=>nx10876, A1=>adderInput_6(14));
   ix10978 : xor2 port map ( Y=>nx10977, A0=>nx10874, A1=>adderInput_6(15));
   ix4935 : xor2 port map ( Y=>label_5(0), A0=>adderInput_5(0), A1=>
      booth_integration_output_5_0);
   ix5662 : mux21_ni port map ( Y=>nx5661, A0=>booth_integration_output_5_0, 
      A1=>nx4778, S0=>nx14482);
   ix4779 : mux21_ni port map ( Y=>nx4778, A0=>neuron(0), A1=>
      booth_integration_output_5_1, S0=>nx14730);
   ix5652 : mux21_ni port map ( Y=>nx5651, A0=>booth_integration_output_5_1, 
      A1=>nx4766, S0=>nx14482);
   ix4767 : mux21_ni port map ( Y=>nx4766, A0=>neuron(1), A1=>
      booth_integration_output_5_2, S0=>nx14730);
   ix5642 : mux21_ni port map ( Y=>nx5641, A0=>booth_integration_output_5_2, 
      A1=>nx4754, S0=>nx14482);
   ix4755 : mux21_ni port map ( Y=>nx4754, A0=>neuron(2), A1=>
      booth_integration_output_5_3, S0=>nx14730);
   ix5632 : mux21_ni port map ( Y=>nx5631, A0=>booth_integration_output_5_3, 
      A1=>nx4742, S0=>nx14482);
   ix4743 : mux21_ni port map ( Y=>nx4742, A0=>neuron(3), A1=>
      booth_integration_output_5_4, S0=>nx14730);
   ix5622 : mux21_ni port map ( Y=>nx5621, A0=>booth_integration_output_5_4, 
      A1=>nx4730, S0=>nx14482);
   ix4731 : mux21_ni port map ( Y=>nx4730, A0=>neuron(4), A1=>
      booth_integration_output_5_5, S0=>nx14730);
   ix5612 : mux21_ni port map ( Y=>nx5611, A0=>booth_integration_output_5_5, 
      A1=>nx4718, S0=>nx14482);
   ix4719 : mux21_ni port map ( Y=>nx4718, A0=>neuron(5), A1=>
      booth_integration_output_5_6, S0=>nx14732);
   ix5602 : mux21_ni port map ( Y=>nx5601, A0=>booth_integration_output_5_6, 
      A1=>nx4706, S0=>nx14482);
   ix4707 : mux21_ni port map ( Y=>nx4706, A0=>neuron(6), A1=>
      booth_integration_output_5_7, S0=>nx14732);
   ix5592 : mux21_ni port map ( Y=>nx5591, A0=>booth_integration_output_5_7, 
      A1=>nx4694, S0=>nx14722);
   ix4695 : mux21_ni port map ( Y=>nx4694, A0=>neuron(7), A1=>
      booth_integration_output_5_8, S0=>nx14732);
   ix5582 : mux21_ni port map ( Y=>nx5581, A0=>booth_integration_output_5_8, 
      A1=>nx4682, S0=>nx14722);
   ix4683 : mux21_ni port map ( Y=>nx4682, A0=>neuron(8), A1=>
      booth_integration_output_5_9, S0=>nx14732);
   ix5572 : mux21_ni port map ( Y=>nx5571, A0=>booth_integration_output_5_9, 
      A1=>nx4670, S0=>nx14722);
   ix4671 : mux21_ni port map ( Y=>nx4670, A0=>neuron(9), A1=>
      booth_integration_output_5_10, S0=>nx14732);
   ix5562 : mux21_ni port map ( Y=>nx5561, A0=>booth_integration_output_5_10, 
      A1=>nx4658, S0=>nx14724);
   ix4659 : mux21_ni port map ( Y=>nx4658, A0=>neuron(10), A1=>
      booth_integration_output_5_11, S0=>nx14732);
   ix5552 : mux21_ni port map ( Y=>nx5551, A0=>booth_integration_output_5_11, 
      A1=>nx4646, S0=>nx14724);
   ix4647 : mux21_ni port map ( Y=>nx4646, A0=>neuron(11), A1=>
      booth_integration_output_5_12, S0=>nx14732);
   ix5542 : mux21_ni port map ( Y=>nx5541, A0=>booth_integration_output_5_12, 
      A1=>nx4634, S0=>nx14724);
   ix4635 : mux21_ni port map ( Y=>nx4634, A0=>neuron(12), A1=>
      booth_integration_output_5_13, S0=>nx14734);
   ix5532 : mux21_ni port map ( Y=>nx5531, A0=>booth_integration_output_5_13, 
      A1=>nx4622, S0=>nx14724);
   ix4623 : mux21_ni port map ( Y=>nx4622, A0=>neuron(13), A1=>
      booth_integration_output_5_14, S0=>nx14734);
   ix5522 : mux21_ni port map ( Y=>nx5521, A0=>booth_integration_output_5_14, 
      A1=>nx4610, S0=>nx14724);
   ix4611 : mux21_ni port map ( Y=>nx4610, A0=>neuron(14), A1=>
      booth_integration_output_5_15, S0=>nx14734);
   ix5512 : mux21 port map ( Y=>nx5511, A0=>nx11397, A1=>nx11028, S0=>
      nx14724);
   ix5162 : mux21_ni port map ( Y=>nx5161, A0=>
      booth_integrtaion_5_shift_Reg_count_0, A1=>nx14262, S0=>nx14628);
   ix5148 : and02 port map ( Y=>nx5147, A0=>nx14838, A1=>
      booth_integrtaion_5_shift_Reg_count_0);
   ix5342 : mux21_ni port map ( Y=>nx5341, A0=>
      booth_integrtaion_5_shift_Reg_count_9, A1=>nx14248, S0=>nx14628);
   ix5332 : mux21_ni port map ( Y=>nx5331, A0=>
      booth_integrtaion_5_shift_Reg_count_9, A1=>
      booth_integrtaion_5_shift_Reg_output_8, S0=>nx14724);
   ix5322 : mux21_ni port map ( Y=>nx5321, A0=>
      booth_integrtaion_5_shift_Reg_count_8, A1=>
      booth_integrtaion_5_shift_Reg_output_8, S0=>nx14628);
   ix5312 : mux21_ni port map ( Y=>nx5311, A0=>
      booth_integrtaion_5_shift_Reg_count_8, A1=>
      booth_integrtaion_5_shift_Reg_output_7, S0=>nx14726);
   ix5302 : mux21_ni port map ( Y=>nx5301, A0=>
      booth_integrtaion_5_shift_Reg_count_7, A1=>
      booth_integrtaion_5_shift_Reg_output_7, S0=>nx14628);
   ix5292 : mux21_ni port map ( Y=>nx5291, A0=>
      booth_integrtaion_5_shift_Reg_count_7, A1=>
      booth_integrtaion_5_shift_Reg_output_6, S0=>nx14726);
   ix5282 : mux21_ni port map ( Y=>nx5281, A0=>
      booth_integrtaion_5_shift_Reg_count_6, A1=>
      booth_integrtaion_5_shift_Reg_output_6, S0=>nx14628);
   ix5272 : mux21_ni port map ( Y=>nx5271, A0=>
      booth_integrtaion_5_shift_Reg_count_6, A1=>
      booth_integrtaion_5_shift_Reg_output_5, S0=>nx14726);
   ix5262 : mux21_ni port map ( Y=>nx5261, A0=>
      booth_integrtaion_5_shift_Reg_count_5, A1=>
      booth_integrtaion_5_shift_Reg_output_5, S0=>nx14628);
   ix5252 : mux21_ni port map ( Y=>nx5251, A0=>
      booth_integrtaion_5_shift_Reg_count_5, A1=>
      booth_integrtaion_5_shift_Reg_output_4, S0=>nx14726);
   ix5242 : mux21_ni port map ( Y=>nx5241, A0=>
      booth_integrtaion_5_shift_Reg_count_4, A1=>
      booth_integrtaion_5_shift_Reg_output_4, S0=>nx14630);
   ix5232 : mux21_ni port map ( Y=>nx5231, A0=>
      booth_integrtaion_5_shift_Reg_count_4, A1=>
      booth_integrtaion_5_shift_Reg_output_3, S0=>nx14726);
   ix5222 : mux21_ni port map ( Y=>nx5221, A0=>
      booth_integrtaion_5_shift_Reg_count_3, A1=>
      booth_integrtaion_5_shift_Reg_output_3, S0=>nx14630);
   ix5212 : mux21_ni port map ( Y=>nx5211, A0=>
      booth_integrtaion_5_shift_Reg_count_3, A1=>
      booth_integrtaion_5_shift_Reg_output_2, S0=>nx14726);
   ix5202 : mux21_ni port map ( Y=>nx5201, A0=>
      booth_integrtaion_5_shift_Reg_count_2, A1=>
      booth_integrtaion_5_shift_Reg_output_2, S0=>nx14630);
   ix5192 : mux21_ni port map ( Y=>nx5191, A0=>
      booth_integrtaion_5_shift_Reg_count_2, A1=>
      booth_integrtaion_5_shift_Reg_output_1, S0=>nx14726);
   ix5182 : mux21_ni port map ( Y=>nx5181, A0=>
      booth_integrtaion_5_shift_Reg_count_1, A1=>
      booth_integrtaion_5_shift_Reg_output_1, S0=>nx14630);
   ix5172 : mux21_ni port map ( Y=>nx5171, A0=>
      booth_integrtaion_5_shift_Reg_count_1, A1=>nx14262, S0=>nx14728);
   ix4051 : and02 port map ( Y=>nx4050, A0=>nx11101, A1=>
      booth_integration_output_5_0);
   ix11104 : or03 port map ( Y=>nx11103, A0=>nx10980, A1=>
      booth_integrtaion_5_shift_reg_output_0, A2=>nx14838);
   ix5502 : mux21_ni port map ( Y=>nx5501, A0=>
      booth_integrtaion_5_booth_output_16, A1=>nx4580, S0=>nx14728);
   ix4581 : nor02ii port map ( Y=>nx4580, A0=>nx11111, A1=>nx14734);
   ix4057 : nor02ii port map ( Y=>nx4056, A0=>nx11096, A1=>
      booth_integrtaion_5_booth_output_16);
   ix4575 : xor2 port map ( Y=>nx2921, A0=>nx11117, A1=>nx11393);
   ix4563 : xor2 port map ( Y=>nx2923, A0=>nx11131, A1=>nx14488);
   ix5472 : mux21_ni port map ( Y=>nx5471, A0=>
      booth_integrtaion_5_booth_output_19, A1=>nx4544, S0=>nx14728);
   ix4545 : nor02ii port map ( Y=>nx4544, A0=>nx11149, A1=>nx14734);
   ix11163 : nor02_2x port map ( Y=>nx4046, A0=>nx11101, A1=>
      booth_integration_output_5_0);
   ix11166 : xor2 port map ( Y=>nx11165, A0=>nx11169, A1=>nx4152);
   ix5452 : mux21_ni port map ( Y=>nx5451, A0=>
      booth_integrtaion_5_booth_output_21, A1=>nx4520, S0=>nx14728);
   ix4521 : nor02ii port map ( Y=>nx4520, A0=>nx11189, A1=>nx14734);
   ix11202 : xor2 port map ( Y=>nx11201, A0=>nx11205, A1=>nx4200);
   ix5432 : mux21_ni port map ( Y=>nx5431, A0=>
      booth_integrtaion_5_booth_output_23, A1=>nx4496, S0=>nx14728);
   ix4497 : nor02ii port map ( Y=>nx4496, A0=>nx11225, A1=>nx14734);
   ix11238 : xor2 port map ( Y=>nx11237, A0=>nx11241, A1=>nx4248);
   ix5412 : mux21_ni port map ( Y=>nx5411, A0=>
      booth_integrtaion_5_booth_output_25, A1=>nx4472, S0=>nx14728);
   ix4473 : nor02ii port map ( Y=>nx4472, A0=>nx11261, A1=>nx14736);
   ix11274 : xor2 port map ( Y=>nx11273, A0=>nx11277, A1=>nx4296);
   ix5392 : mux21_ni port map ( Y=>nx5391, A0=>
      booth_integrtaion_5_booth_output_27, A1=>nx4448, S0=>nx14728);
   ix4449 : nor02ii port map ( Y=>nx4448, A0=>nx11297, A1=>nx14736);
   ix11310 : xor2 port map ( Y=>nx11309, A0=>nx11313, A1=>nx4344);
   ix5372 : mux21_ni port map ( Y=>nx5371, A0=>
      booth_integrtaion_5_booth_output_29, A1=>nx4424, S0=>nx14480);
   ix4425 : nor02ii port map ( Y=>nx4424, A0=>nx11333, A1=>nx14736);
   ix11346 : xor2 port map ( Y=>nx11345, A0=>nx11353, A1=>nx4392);
   ix5362 : mux21_ni port map ( Y=>nx5361, A0=>
      booth_integrtaion_5_booth_output_31, A1=>nx4412, S0=>nx14480);
   ix4413 : nor02ii port map ( Y=>nx4412, A0=>nx11350, A1=>nx14736);
   ix4407 : xor2 port map ( Y=>nx4406, A0=>nx11353, A1=>nx11365);
   ix4593 : nor02ii port map ( Y=>nx4592, A0=>nx4056, A1=>nx14736);
   ix11423 : xor2 port map ( Y=>nx11422, A0=>nx11411, A1=>adderInput_5(2));
   ix11435 : xor2 port map ( Y=>nx11434, A0=>nx11409, A1=>adderInput_5(4));
   ix11447 : xor2 port map ( Y=>nx11446, A0=>nx11407, A1=>adderInput_5(6));
   ix11459 : xor2 port map ( Y=>nx11458, A0=>nx11405, A1=>adderInput_5(8));
   ix11471 : xor2 port map ( Y=>nx11470, A0=>nx11403, A1=>adderInput_5(10));
   ix11483 : xor2 port map ( Y=>nx11482, A0=>nx11401, A1=>adderInput_5(12));
   ix11495 : xor2 port map ( Y=>nx11494, A0=>nx11399, A1=>adderInput_5(14));
   ix11501 : xor2 port map ( Y=>nx11500, A0=>nx11397, A1=>adderInput_5(15));
   ix5921 : xor2 port map ( Y=>label_4(0), A0=>adderInput_4(0), A1=>
      booth_integration_output_4_0);
   ix6192 : mux21_ni port map ( Y=>nx6191, A0=>booth_integration_output_4_0, 
      A1=>nx5764, S0=>nx14504);
   ix5765 : mux21_ni port map ( Y=>nx5764, A0=>neuron(0), A1=>
      booth_integration_output_4_1, S0=>nx14746);
   ix6182 : mux21_ni port map ( Y=>nx6181, A0=>booth_integration_output_4_1, 
      A1=>nx5752, S0=>nx14504);
   ix5753 : mux21_ni port map ( Y=>nx5752, A0=>neuron(1), A1=>
      booth_integration_output_4_2, S0=>nx14746);
   ix6172 : mux21_ni port map ( Y=>nx6171, A0=>booth_integration_output_4_2, 
      A1=>nx5740, S0=>nx14504);
   ix5741 : mux21_ni port map ( Y=>nx5740, A0=>neuron(2), A1=>
      booth_integration_output_4_3, S0=>nx14746);
   ix6162 : mux21_ni port map ( Y=>nx6161, A0=>booth_integration_output_4_3, 
      A1=>nx5728, S0=>nx14504);
   ix5729 : mux21_ni port map ( Y=>nx5728, A0=>neuron(3), A1=>
      booth_integration_output_4_4, S0=>nx14746);
   ix6152 : mux21_ni port map ( Y=>nx6151, A0=>booth_integration_output_4_4, 
      A1=>nx5716, S0=>nx14504);
   ix5717 : mux21_ni port map ( Y=>nx5716, A0=>neuron(4), A1=>
      booth_integration_output_4_5, S0=>nx14746);
   ix6142 : mux21_ni port map ( Y=>nx6141, A0=>booth_integration_output_4_5, 
      A1=>nx5704, S0=>nx14504);
   ix5705 : mux21_ni port map ( Y=>nx5704, A0=>neuron(5), A1=>
      booth_integration_output_4_6, S0=>nx14748);
   ix6132 : mux21_ni port map ( Y=>nx6131, A0=>booth_integration_output_4_6, 
      A1=>nx5692, S0=>nx14504);
   ix5693 : mux21_ni port map ( Y=>nx5692, A0=>neuron(6), A1=>
      booth_integration_output_4_7, S0=>nx14748);
   ix6122 : mux21_ni port map ( Y=>nx6121, A0=>booth_integration_output_4_7, 
      A1=>nx5680, S0=>nx14738);
   ix5681 : mux21_ni port map ( Y=>nx5680, A0=>neuron(7), A1=>
      booth_integration_output_4_8, S0=>nx14748);
   ix6112 : mux21_ni port map ( Y=>nx6111, A0=>booth_integration_output_4_8, 
      A1=>nx5668, S0=>nx14738);
   ix5669 : mux21_ni port map ( Y=>nx5668, A0=>neuron(8), A1=>
      booth_integration_output_4_9, S0=>nx14748);
   ix6102 : mux21_ni port map ( Y=>nx6101, A0=>booth_integration_output_4_9, 
      A1=>nx5656, S0=>nx14738);
   ix5657 : mux21_ni port map ( Y=>nx5656, A0=>neuron(9), A1=>
      booth_integration_output_4_10, S0=>nx14748);
   ix6092 : mux21_ni port map ( Y=>nx6091, A0=>booth_integration_output_4_10, 
      A1=>nx5644, S0=>nx14740);
   ix5645 : mux21_ni port map ( Y=>nx5644, A0=>neuron(10), A1=>
      booth_integration_output_4_11, S0=>nx14748);
   ix6082 : mux21_ni port map ( Y=>nx6081, A0=>booth_integration_output_4_11, 
      A1=>nx5632, S0=>nx14740);
   ix5633 : mux21_ni port map ( Y=>nx5632, A0=>neuron(11), A1=>
      booth_integration_output_4_12, S0=>nx14748);
   ix6072 : mux21_ni port map ( Y=>nx6071, A0=>booth_integration_output_4_12, 
      A1=>nx5620, S0=>nx14740);
   ix5621 : mux21_ni port map ( Y=>nx5620, A0=>neuron(12), A1=>
      booth_integration_output_4_13, S0=>nx14750);
   ix6062 : mux21_ni port map ( Y=>nx6061, A0=>booth_integration_output_4_13, 
      A1=>nx5608, S0=>nx14740);
   ix5609 : mux21_ni port map ( Y=>nx5608, A0=>neuron(13), A1=>
      booth_integration_output_4_14, S0=>nx14750);
   ix6052 : mux21_ni port map ( Y=>nx6051, A0=>booth_integration_output_4_14, 
      A1=>nx5596, S0=>nx14740);
   ix5597 : mux21_ni port map ( Y=>nx5596, A0=>neuron(14), A1=>
      booth_integration_output_4_15, S0=>nx14750);
   ix6042 : mux21 port map ( Y=>nx6041, A0=>nx11920, A1=>nx11551, S0=>
      nx14740);
   ix5692 : mux21_ni port map ( Y=>nx5691, A0=>
      booth_integrtaion_4_shift_Reg_count_0, A1=>nx14284, S0=>nx14632);
   ix5678 : and02 port map ( Y=>nx5677, A0=>nx14842, A1=>
      booth_integrtaion_4_shift_Reg_count_0);
   ix5872 : mux21_ni port map ( Y=>nx5871, A0=>
      booth_integrtaion_4_shift_Reg_count_9, A1=>nx14270, S0=>nx14632);
   ix5862 : mux21_ni port map ( Y=>nx5861, A0=>
      booth_integrtaion_4_shift_Reg_count_9, A1=>
      booth_integrtaion_4_shift_Reg_output_8, S0=>nx14740);
   ix5852 : mux21_ni port map ( Y=>nx5851, A0=>
      booth_integrtaion_4_shift_Reg_count_8, A1=>
      booth_integrtaion_4_shift_Reg_output_8, S0=>nx14632);
   ix5842 : mux21_ni port map ( Y=>nx5841, A0=>
      booth_integrtaion_4_shift_Reg_count_8, A1=>
      booth_integrtaion_4_shift_Reg_output_7, S0=>nx14742);
   ix5832 : mux21_ni port map ( Y=>nx5831, A0=>
      booth_integrtaion_4_shift_Reg_count_7, A1=>
      booth_integrtaion_4_shift_Reg_output_7, S0=>nx14632);
   ix5822 : mux21_ni port map ( Y=>nx5821, A0=>
      booth_integrtaion_4_shift_Reg_count_7, A1=>
      booth_integrtaion_4_shift_Reg_output_6, S0=>nx14742);
   ix5812 : mux21_ni port map ( Y=>nx5811, A0=>
      booth_integrtaion_4_shift_Reg_count_6, A1=>
      booth_integrtaion_4_shift_Reg_output_6, S0=>nx14632);
   ix5802 : mux21_ni port map ( Y=>nx5801, A0=>
      booth_integrtaion_4_shift_Reg_count_6, A1=>
      booth_integrtaion_4_shift_Reg_output_5, S0=>nx14742);
   ix5792 : mux21_ni port map ( Y=>nx5791, A0=>
      booth_integrtaion_4_shift_Reg_count_5, A1=>
      booth_integrtaion_4_shift_Reg_output_5, S0=>nx14632);
   ix5782 : mux21_ni port map ( Y=>nx5781, A0=>
      booth_integrtaion_4_shift_Reg_count_5, A1=>
      booth_integrtaion_4_shift_Reg_output_4, S0=>nx14742);
   ix5772 : mux21_ni port map ( Y=>nx5771, A0=>
      booth_integrtaion_4_shift_Reg_count_4, A1=>
      booth_integrtaion_4_shift_Reg_output_4, S0=>nx14634);
   ix5762 : mux21_ni port map ( Y=>nx5761, A0=>
      booth_integrtaion_4_shift_Reg_count_4, A1=>
      booth_integrtaion_4_shift_Reg_output_3, S0=>nx14742);
   ix5752 : mux21_ni port map ( Y=>nx5751, A0=>
      booth_integrtaion_4_shift_Reg_count_3, A1=>
      booth_integrtaion_4_shift_Reg_output_3, S0=>nx14634);
   ix5742 : mux21_ni port map ( Y=>nx5741, A0=>
      booth_integrtaion_4_shift_Reg_count_3, A1=>
      booth_integrtaion_4_shift_Reg_output_2, S0=>nx14742);
   ix5732 : mux21_ni port map ( Y=>nx5731, A0=>
      booth_integrtaion_4_shift_Reg_count_2, A1=>
      booth_integrtaion_4_shift_Reg_output_2, S0=>nx14634);
   ix5722 : mux21_ni port map ( Y=>nx5721, A0=>
      booth_integrtaion_4_shift_Reg_count_2, A1=>
      booth_integrtaion_4_shift_Reg_output_1, S0=>nx14742);
   ix5712 : mux21_ni port map ( Y=>nx5711, A0=>
      booth_integrtaion_4_shift_Reg_count_1, A1=>
      booth_integrtaion_4_shift_Reg_output_1, S0=>nx14634);
   ix5702 : mux21_ni port map ( Y=>nx5701, A0=>
      booth_integrtaion_4_shift_Reg_count_1, A1=>nx14284, S0=>nx14744);
   ix5037 : and02 port map ( Y=>nx5036, A0=>nx11624, A1=>
      booth_integration_output_4_0);
   ix11627 : or03 port map ( Y=>nx11626, A0=>nx11503, A1=>
      booth_integrtaion_4_shift_reg_output_0, A2=>nx14842);
   ix6032 : mux21_ni port map ( Y=>nx6031, A0=>
      booth_integrtaion_4_booth_output_16, A1=>nx5566, S0=>nx14744);
   ix5567 : nor02ii port map ( Y=>nx5566, A0=>nx11634, A1=>nx14750);
   ix5043 : nor02ii port map ( Y=>nx5042, A0=>nx11619, A1=>
      booth_integrtaion_4_booth_output_16);
   ix5561 : xor2 port map ( Y=>nx2939, A0=>nx11640, A1=>nx11916);
   ix5549 : xor2 port map ( Y=>nx2940, A0=>nx11654, A1=>nx14510);
   ix6002 : mux21_ni port map ( Y=>nx6001, A0=>
      booth_integrtaion_4_booth_output_19, A1=>nx5530, S0=>nx14744);
   ix5531 : nor02ii port map ( Y=>nx5530, A0=>nx11672, A1=>nx14750);
   ix11686 : nor02_2x port map ( Y=>nx5032, A0=>nx11624, A1=>
      booth_integration_output_4_0);
   ix11689 : xor2 port map ( Y=>nx11688, A0=>nx11692, A1=>nx5138);
   ix5982 : mux21_ni port map ( Y=>nx5981, A0=>
      booth_integrtaion_4_booth_output_21, A1=>nx5506, S0=>nx14744);
   ix5507 : nor02ii port map ( Y=>nx5506, A0=>nx11712, A1=>nx14750);
   ix11725 : xor2 port map ( Y=>nx11724, A0=>nx11728, A1=>nx5186);
   ix5962 : mux21_ni port map ( Y=>nx5961, A0=>
      booth_integrtaion_4_booth_output_23, A1=>nx5482, S0=>nx14744);
   ix5483 : nor02ii port map ( Y=>nx5482, A0=>nx11748, A1=>nx14750);
   ix11761 : xor2 port map ( Y=>nx11760, A0=>nx11764, A1=>nx5234);
   ix5942 : mux21_ni port map ( Y=>nx5941, A0=>
      booth_integrtaion_4_booth_output_25, A1=>nx5458, S0=>nx14744);
   ix5459 : nor02ii port map ( Y=>nx5458, A0=>nx11784, A1=>nx14752);
   ix11797 : xor2 port map ( Y=>nx11796, A0=>nx11800, A1=>nx5282);
   ix5922 : mux21_ni port map ( Y=>nx5921, A0=>
      booth_integrtaion_4_booth_output_27, A1=>nx5434, S0=>nx14744);
   ix5435 : nor02ii port map ( Y=>nx5434, A0=>nx11820, A1=>nx14752);
   ix11833 : xor2 port map ( Y=>nx11832, A0=>nx11836, A1=>nx5330);
   ix5902 : mux21_ni port map ( Y=>nx5901, A0=>
      booth_integrtaion_4_booth_output_29, A1=>nx5410, S0=>nx14502);
   ix5411 : nor02ii port map ( Y=>nx5410, A0=>nx11856, A1=>nx14752);
   ix11869 : xor2 port map ( Y=>nx11868, A0=>nx11876, A1=>nx5378);
   ix5892 : mux21_ni port map ( Y=>nx5891, A0=>
      booth_integrtaion_4_booth_output_31, A1=>nx5398, S0=>nx14502);
   ix5399 : nor02ii port map ( Y=>nx5398, A0=>nx11873, A1=>nx14752);
   ix5393 : xor2 port map ( Y=>nx5392, A0=>nx11876, A1=>nx11888);
   ix5579 : nor02ii port map ( Y=>nx5578, A0=>nx5042, A1=>nx14752);
   ix11946 : xor2 port map ( Y=>nx11945, A0=>nx11934, A1=>adderInput_4(2));
   ix11958 : xor2 port map ( Y=>nx11957, A0=>nx11932, A1=>adderInput_4(4));
   ix11970 : xor2 port map ( Y=>nx11969, A0=>nx11930, A1=>adderInput_4(6));
   ix11982 : xor2 port map ( Y=>nx11981, A0=>nx11928, A1=>adderInput_4(8));
   ix11994 : xor2 port map ( Y=>nx11993, A0=>nx11926, A1=>adderInput_4(10));
   ix12006 : xor2 port map ( Y=>nx12005, A0=>nx11924, A1=>adderInput_4(12));
   ix12018 : xor2 port map ( Y=>nx12017, A0=>nx11922, A1=>adderInput_4(14));
   ix12024 : xor2 port map ( Y=>nx12023, A0=>nx11920, A1=>adderInput_4(15));
   ix6907 : xor2 port map ( Y=>label_3(0), A0=>adderInput_3(0), A1=>
      booth_integration_output_3_0);
   ix6722 : mux21_ni port map ( Y=>nx6721, A0=>booth_integration_output_3_0, 
      A1=>nx6750, S0=>nx14526);
   ix6751 : mux21_ni port map ( Y=>nx6750, A0=>neuron(0), A1=>
      booth_integration_output_3_1, S0=>nx14762);
   ix6712 : mux21_ni port map ( Y=>nx6711, A0=>booth_integration_output_3_1, 
      A1=>nx6738, S0=>nx14526);
   ix6739 : mux21_ni port map ( Y=>nx6738, A0=>neuron(1), A1=>
      booth_integration_output_3_2, S0=>nx14762);
   ix6702 : mux21_ni port map ( Y=>nx6701, A0=>booth_integration_output_3_2, 
      A1=>nx6726, S0=>nx14526);
   ix6727 : mux21_ni port map ( Y=>nx6726, A0=>neuron(2), A1=>
      booth_integration_output_3_3, S0=>nx14762);
   ix6692 : mux21_ni port map ( Y=>nx6691, A0=>booth_integration_output_3_3, 
      A1=>nx6714, S0=>nx14526);
   ix6715 : mux21_ni port map ( Y=>nx6714, A0=>neuron(3), A1=>
      booth_integration_output_3_4, S0=>nx14762);
   ix6682 : mux21_ni port map ( Y=>nx6681, A0=>booth_integration_output_3_4, 
      A1=>nx6702, S0=>nx14526);
   ix6703 : mux21_ni port map ( Y=>nx6702, A0=>neuron(4), A1=>
      booth_integration_output_3_5, S0=>nx14762);
   ix6672 : mux21_ni port map ( Y=>nx6671, A0=>booth_integration_output_3_5, 
      A1=>nx6690, S0=>nx14526);
   ix6691 : mux21_ni port map ( Y=>nx6690, A0=>neuron(5), A1=>
      booth_integration_output_3_6, S0=>nx14764);
   ix6662 : mux21_ni port map ( Y=>nx6661, A0=>booth_integration_output_3_6, 
      A1=>nx6678, S0=>nx14526);
   ix6679 : mux21_ni port map ( Y=>nx6678, A0=>neuron(6), A1=>
      booth_integration_output_3_7, S0=>nx14764);
   ix6652 : mux21_ni port map ( Y=>nx6651, A0=>booth_integration_output_3_7, 
      A1=>nx6666, S0=>nx14754);
   ix6667 : mux21_ni port map ( Y=>nx6666, A0=>neuron(7), A1=>
      booth_integration_output_3_8, S0=>nx14764);
   ix6642 : mux21_ni port map ( Y=>nx6641, A0=>booth_integration_output_3_8, 
      A1=>nx6654, S0=>nx14754);
   ix6655 : mux21_ni port map ( Y=>nx6654, A0=>neuron(8), A1=>
      booth_integration_output_3_9, S0=>nx14764);
   ix6632 : mux21_ni port map ( Y=>nx6631, A0=>booth_integration_output_3_9, 
      A1=>nx6642, S0=>nx14754);
   ix6643 : mux21_ni port map ( Y=>nx6642, A0=>neuron(9), A1=>
      booth_integration_output_3_10, S0=>nx14764);
   ix6622 : mux21_ni port map ( Y=>nx6621, A0=>booth_integration_output_3_10, 
      A1=>nx6630, S0=>nx14756);
   ix6631 : mux21_ni port map ( Y=>nx6630, A0=>neuron(10), A1=>
      booth_integration_output_3_11, S0=>nx14764);
   ix6612 : mux21_ni port map ( Y=>nx6611, A0=>booth_integration_output_3_11, 
      A1=>nx6618, S0=>nx14756);
   ix6619 : mux21_ni port map ( Y=>nx6618, A0=>neuron(11), A1=>
      booth_integration_output_3_12, S0=>nx14764);
   ix6602 : mux21_ni port map ( Y=>nx6601, A0=>booth_integration_output_3_12, 
      A1=>nx6606, S0=>nx14756);
   ix6607 : mux21_ni port map ( Y=>nx6606, A0=>neuron(12), A1=>
      booth_integration_output_3_13, S0=>nx14766);
   ix6592 : mux21_ni port map ( Y=>nx6591, A0=>booth_integration_output_3_13, 
      A1=>nx6594, S0=>nx14756);
   ix6595 : mux21_ni port map ( Y=>nx6594, A0=>neuron(13), A1=>
      booth_integration_output_3_14, S0=>nx14766);
   ix6582 : mux21_ni port map ( Y=>nx6581, A0=>booth_integration_output_3_14, 
      A1=>nx6582, S0=>nx14756);
   ix6583 : mux21_ni port map ( Y=>nx6582, A0=>neuron(14), A1=>
      booth_integration_output_3_15, S0=>nx14766);
   ix6572 : mux21 port map ( Y=>nx6571, A0=>nx12443, A1=>nx12074, S0=>
      nx14756);
   ix6222 : mux21_ni port map ( Y=>nx6221, A0=>
      booth_integrtaion_3_shift_Reg_count_0, A1=>nx14306, S0=>nx14636);
   ix6208 : and02 port map ( Y=>nx6207, A0=>nx14846, A1=>
      booth_integrtaion_3_shift_Reg_count_0);
   ix6402 : mux21_ni port map ( Y=>nx6401, A0=>
      booth_integrtaion_3_shift_Reg_count_9, A1=>nx14292, S0=>nx14636);
   ix6392 : mux21_ni port map ( Y=>nx6391, A0=>
      booth_integrtaion_3_shift_Reg_count_9, A1=>
      booth_integrtaion_3_shift_Reg_output_8, S0=>nx14756);
   ix6382 : mux21_ni port map ( Y=>nx6381, A0=>
      booth_integrtaion_3_shift_Reg_count_8, A1=>
      booth_integrtaion_3_shift_Reg_output_8, S0=>nx14636);
   ix6372 : mux21_ni port map ( Y=>nx6371, A0=>
      booth_integrtaion_3_shift_Reg_count_8, A1=>
      booth_integrtaion_3_shift_Reg_output_7, S0=>nx14758);
   ix6362 : mux21_ni port map ( Y=>nx6361, A0=>
      booth_integrtaion_3_shift_Reg_count_7, A1=>
      booth_integrtaion_3_shift_Reg_output_7, S0=>nx14636);
   ix6352 : mux21_ni port map ( Y=>nx6351, A0=>
      booth_integrtaion_3_shift_Reg_count_7, A1=>
      booth_integrtaion_3_shift_Reg_output_6, S0=>nx14758);
   ix6342 : mux21_ni port map ( Y=>nx6341, A0=>
      booth_integrtaion_3_shift_Reg_count_6, A1=>
      booth_integrtaion_3_shift_Reg_output_6, S0=>nx14636);
   ix6332 : mux21_ni port map ( Y=>nx6331, A0=>
      booth_integrtaion_3_shift_Reg_count_6, A1=>
      booth_integrtaion_3_shift_Reg_output_5, S0=>nx14758);
   ix6322 : mux21_ni port map ( Y=>nx6321, A0=>
      booth_integrtaion_3_shift_Reg_count_5, A1=>
      booth_integrtaion_3_shift_Reg_output_5, S0=>nx14636);
   ix6312 : mux21_ni port map ( Y=>nx6311, A0=>
      booth_integrtaion_3_shift_Reg_count_5, A1=>
      booth_integrtaion_3_shift_Reg_output_4, S0=>nx14758);
   ix6302 : mux21_ni port map ( Y=>nx6301, A0=>
      booth_integrtaion_3_shift_Reg_count_4, A1=>
      booth_integrtaion_3_shift_Reg_output_4, S0=>nx14638);
   ix6292 : mux21_ni port map ( Y=>nx6291, A0=>
      booth_integrtaion_3_shift_Reg_count_4, A1=>
      booth_integrtaion_3_shift_Reg_output_3, S0=>nx14758);
   ix6282 : mux21_ni port map ( Y=>nx6281, A0=>
      booth_integrtaion_3_shift_Reg_count_3, A1=>
      booth_integrtaion_3_shift_Reg_output_3, S0=>nx14638);
   ix6272 : mux21_ni port map ( Y=>nx6271, A0=>
      booth_integrtaion_3_shift_Reg_count_3, A1=>
      booth_integrtaion_3_shift_Reg_output_2, S0=>nx14758);
   ix6262 : mux21_ni port map ( Y=>nx6261, A0=>
      booth_integrtaion_3_shift_Reg_count_2, A1=>
      booth_integrtaion_3_shift_Reg_output_2, S0=>nx14638);
   ix6252 : mux21_ni port map ( Y=>nx6251, A0=>
      booth_integrtaion_3_shift_Reg_count_2, A1=>
      booth_integrtaion_3_shift_Reg_output_1, S0=>nx14758);
   ix6242 : mux21_ni port map ( Y=>nx6241, A0=>
      booth_integrtaion_3_shift_Reg_count_1, A1=>
      booth_integrtaion_3_shift_Reg_output_1, S0=>nx14638);
   ix6232 : mux21_ni port map ( Y=>nx6231, A0=>
      booth_integrtaion_3_shift_Reg_count_1, A1=>nx14306, S0=>nx14760);
   ix6023 : and02 port map ( Y=>nx6022, A0=>nx12147, A1=>
      booth_integration_output_3_0);
   ix12150 : or03 port map ( Y=>nx12149, A0=>nx12026, A1=>
      booth_integrtaion_3_shift_reg_output_0, A2=>nx14846);
   ix6562 : mux21_ni port map ( Y=>nx6561, A0=>
      booth_integrtaion_3_booth_output_16, A1=>nx6552, S0=>nx14760);
   ix6553 : nor02ii port map ( Y=>nx6552, A0=>nx12157, A1=>nx14766);
   ix6029 : nor02ii port map ( Y=>nx6028, A0=>nx12142, A1=>
      booth_integrtaion_3_booth_output_16);
   ix6547 : xor2 port map ( Y=>nx2954, A0=>nx12163, A1=>nx12439);
   ix6535 : xor2 port map ( Y=>nx2955, A0=>nx12177, A1=>nx14532);
   ix6532 : mux21_ni port map ( Y=>nx6531, A0=>
      booth_integrtaion_3_booth_output_19, A1=>nx6516, S0=>nx14760);
   ix6517 : nor02ii port map ( Y=>nx6516, A0=>nx12195, A1=>nx14766);
   ix12209 : nor02_2x port map ( Y=>nx6018, A0=>nx12147, A1=>
      booth_integration_output_3_0);
   ix12212 : xor2 port map ( Y=>nx12211, A0=>nx12215, A1=>nx6124);
   ix6512 : mux21_ni port map ( Y=>nx6511, A0=>
      booth_integrtaion_3_booth_output_21, A1=>nx6492, S0=>nx14760);
   ix6493 : nor02ii port map ( Y=>nx6492, A0=>nx12235, A1=>nx14766);
   ix12248 : xor2 port map ( Y=>nx12247, A0=>nx12251, A1=>nx6172);
   ix6492 : mux21_ni port map ( Y=>nx6491, A0=>
      booth_integrtaion_3_booth_output_23, A1=>nx6468, S0=>nx14760);
   ix6469 : nor02ii port map ( Y=>nx6468, A0=>nx12271, A1=>nx14766);
   ix12284 : xor2 port map ( Y=>nx12283, A0=>nx12287, A1=>nx6220);
   ix6472 : mux21_ni port map ( Y=>nx6471, A0=>
      booth_integrtaion_3_booth_output_25, A1=>nx6444, S0=>nx14760);
   ix6445 : nor02ii port map ( Y=>nx6444, A0=>nx12307, A1=>nx14768);
   ix12320 : xor2 port map ( Y=>nx12319, A0=>nx12323, A1=>nx6268);
   ix6452 : mux21_ni port map ( Y=>nx6451, A0=>
      booth_integrtaion_3_booth_output_27, A1=>nx6420, S0=>nx14760);
   ix6421 : nor02ii port map ( Y=>nx6420, A0=>nx12343, A1=>nx14768);
   ix12356 : xor2 port map ( Y=>nx12355, A0=>nx12359, A1=>nx6316);
   ix6432 : mux21_ni port map ( Y=>nx6431, A0=>
      booth_integrtaion_3_booth_output_29, A1=>nx6396, S0=>nx14524);
   ix6397 : nor02ii port map ( Y=>nx6396, A0=>nx12379, A1=>nx14768);
   ix12392 : xor2 port map ( Y=>nx12391, A0=>nx12399, A1=>nx6364);
   ix6422 : mux21_ni port map ( Y=>nx6421, A0=>
      booth_integrtaion_3_booth_output_31, A1=>nx6384, S0=>nx14524);
   ix6385 : nor02ii port map ( Y=>nx6384, A0=>nx12396, A1=>nx14768);
   ix6379 : xor2 port map ( Y=>nx6378, A0=>nx12399, A1=>nx12411);
   ix6565 : nor02ii port map ( Y=>nx6564, A0=>nx6028, A1=>nx14768);
   ix12469 : xor2 port map ( Y=>nx12468, A0=>nx12457, A1=>adderInput_3(2));
   ix12481 : xor2 port map ( Y=>nx12480, A0=>nx12455, A1=>adderInput_3(4));
   ix12493 : xor2 port map ( Y=>nx12492, A0=>nx12453, A1=>adderInput_3(6));
   ix12505 : xor2 port map ( Y=>nx12504, A0=>nx12451, A1=>adderInput_3(8));
   ix12517 : xor2 port map ( Y=>nx12516, A0=>nx12449, A1=>adderInput_3(10));
   ix12529 : xor2 port map ( Y=>nx12528, A0=>nx12447, A1=>adderInput_3(12));
   ix12541 : xor2 port map ( Y=>nx12540, A0=>nx12445, A1=>adderInput_3(14));
   ix12547 : xor2 port map ( Y=>nx12546, A0=>nx12443, A1=>adderInput_3(15));
   ix7893 : xor2 port map ( Y=>label_2(0), A0=>adderInput_2(0), A1=>
      booth_integration_output_2_0);
   ix7252 : mux21_ni port map ( Y=>nx7251, A0=>booth_integration_output_2_0, 
      A1=>nx7736, S0=>nx14548);
   ix7737 : mux21_ni port map ( Y=>nx7736, A0=>neuron(0), A1=>
      booth_integration_output_2_1, S0=>nx14778);
   ix7242 : mux21_ni port map ( Y=>nx7241, A0=>booth_integration_output_2_1, 
      A1=>nx7724, S0=>nx14548);
   ix7725 : mux21_ni port map ( Y=>nx7724, A0=>neuron(1), A1=>
      booth_integration_output_2_2, S0=>nx14778);
   ix7232 : mux21_ni port map ( Y=>nx7231, A0=>booth_integration_output_2_2, 
      A1=>nx7712, S0=>nx14548);
   ix7713 : mux21_ni port map ( Y=>nx7712, A0=>neuron(2), A1=>
      booth_integration_output_2_3, S0=>nx14778);
   ix7222 : mux21_ni port map ( Y=>nx7221, A0=>booth_integration_output_2_3, 
      A1=>nx7700, S0=>nx14548);
   ix7701 : mux21_ni port map ( Y=>nx7700, A0=>neuron(3), A1=>
      booth_integration_output_2_4, S0=>nx14778);
   ix7212 : mux21_ni port map ( Y=>nx7211, A0=>booth_integration_output_2_4, 
      A1=>nx7688, S0=>nx14548);
   ix7689 : mux21_ni port map ( Y=>nx7688, A0=>neuron(4), A1=>
      booth_integration_output_2_5, S0=>nx14778);
   ix7202 : mux21_ni port map ( Y=>nx7201, A0=>booth_integration_output_2_5, 
      A1=>nx7676, S0=>nx14548);
   ix7677 : mux21_ni port map ( Y=>nx7676, A0=>neuron(5), A1=>
      booth_integration_output_2_6, S0=>nx14780);
   ix7192 : mux21_ni port map ( Y=>nx7191, A0=>booth_integration_output_2_6, 
      A1=>nx7664, S0=>nx14548);
   ix7665 : mux21_ni port map ( Y=>nx7664, A0=>neuron(6), A1=>
      booth_integration_output_2_7, S0=>nx14780);
   ix7182 : mux21_ni port map ( Y=>nx7181, A0=>booth_integration_output_2_7, 
      A1=>nx7652, S0=>nx14770);
   ix7653 : mux21_ni port map ( Y=>nx7652, A0=>neuron(7), A1=>
      booth_integration_output_2_8, S0=>nx14780);
   ix7172 : mux21_ni port map ( Y=>nx7171, A0=>booth_integration_output_2_8, 
      A1=>nx7640, S0=>nx14770);
   ix7641 : mux21_ni port map ( Y=>nx7640, A0=>neuron(8), A1=>
      booth_integration_output_2_9, S0=>nx14780);
   ix7162 : mux21_ni port map ( Y=>nx7161, A0=>booth_integration_output_2_9, 
      A1=>nx7628, S0=>nx14770);
   ix7629 : mux21_ni port map ( Y=>nx7628, A0=>neuron(9), A1=>
      booth_integration_output_2_10, S0=>nx14780);
   ix7152 : mux21_ni port map ( Y=>nx7151, A0=>booth_integration_output_2_10, 
      A1=>nx7616, S0=>nx14772);
   ix7617 : mux21_ni port map ( Y=>nx7616, A0=>neuron(10), A1=>
      booth_integration_output_2_11, S0=>nx14780);
   ix7142 : mux21_ni port map ( Y=>nx7141, A0=>booth_integration_output_2_11, 
      A1=>nx7604, S0=>nx14772);
   ix7605 : mux21_ni port map ( Y=>nx7604, A0=>neuron(11), A1=>
      booth_integration_output_2_12, S0=>nx14780);
   ix7132 : mux21_ni port map ( Y=>nx7131, A0=>booth_integration_output_2_12, 
      A1=>nx7592, S0=>nx14772);
   ix7593 : mux21_ni port map ( Y=>nx7592, A0=>neuron(12), A1=>
      booth_integration_output_2_13, S0=>nx14782);
   ix7122 : mux21_ni port map ( Y=>nx7121, A0=>booth_integration_output_2_13, 
      A1=>nx7580, S0=>nx14772);
   ix7581 : mux21_ni port map ( Y=>nx7580, A0=>neuron(13), A1=>
      booth_integration_output_2_14, S0=>nx14782);
   ix7112 : mux21_ni port map ( Y=>nx7111, A0=>booth_integration_output_2_14, 
      A1=>nx7568, S0=>nx14772);
   ix7569 : mux21_ni port map ( Y=>nx7568, A0=>neuron(14), A1=>
      booth_integration_output_2_15, S0=>nx14782);
   ix7102 : mux21 port map ( Y=>nx7101, A0=>nx12966, A1=>nx12597, S0=>
      nx14772);
   ix6752 : mux21_ni port map ( Y=>nx6751, A0=>
      booth_integrtaion_2_shift_Reg_count_0, A1=>nx14328, S0=>nx14640);
   ix6738 : and02 port map ( Y=>nx6737, A0=>nx14850, A1=>
      booth_integrtaion_2_shift_Reg_count_0);
   ix6932 : mux21_ni port map ( Y=>nx6931, A0=>
      booth_integrtaion_2_shift_Reg_count_9, A1=>nx14314, S0=>nx14640);
   ix6922 : mux21_ni port map ( Y=>nx6921, A0=>
      booth_integrtaion_2_shift_Reg_count_9, A1=>
      booth_integrtaion_2_shift_Reg_output_8, S0=>nx14772);
   ix6912 : mux21_ni port map ( Y=>nx6911, A0=>
      booth_integrtaion_2_shift_Reg_count_8, A1=>
      booth_integrtaion_2_shift_Reg_output_8, S0=>nx14640);
   ix6902 : mux21_ni port map ( Y=>nx6901, A0=>
      booth_integrtaion_2_shift_Reg_count_8, A1=>
      booth_integrtaion_2_shift_Reg_output_7, S0=>nx14774);
   ix6892 : mux21_ni port map ( Y=>nx6891, A0=>
      booth_integrtaion_2_shift_Reg_count_7, A1=>
      booth_integrtaion_2_shift_Reg_output_7, S0=>nx14640);
   ix6882 : mux21_ni port map ( Y=>nx6881, A0=>
      booth_integrtaion_2_shift_Reg_count_7, A1=>
      booth_integrtaion_2_shift_Reg_output_6, S0=>nx14774);
   ix6872 : mux21_ni port map ( Y=>nx6871, A0=>
      booth_integrtaion_2_shift_Reg_count_6, A1=>
      booth_integrtaion_2_shift_Reg_output_6, S0=>nx14640);
   ix6862 : mux21_ni port map ( Y=>nx6861, A0=>
      booth_integrtaion_2_shift_Reg_count_6, A1=>
      booth_integrtaion_2_shift_Reg_output_5, S0=>nx14774);
   ix6852 : mux21_ni port map ( Y=>nx6851, A0=>
      booth_integrtaion_2_shift_Reg_count_5, A1=>
      booth_integrtaion_2_shift_Reg_output_5, S0=>nx14640);
   ix6842 : mux21_ni port map ( Y=>nx6841, A0=>
      booth_integrtaion_2_shift_Reg_count_5, A1=>
      booth_integrtaion_2_shift_Reg_output_4, S0=>nx14774);
   ix6832 : mux21_ni port map ( Y=>nx6831, A0=>
      booth_integrtaion_2_shift_Reg_count_4, A1=>
      booth_integrtaion_2_shift_Reg_output_4, S0=>nx14642);
   ix6822 : mux21_ni port map ( Y=>nx6821, A0=>
      booth_integrtaion_2_shift_Reg_count_4, A1=>
      booth_integrtaion_2_shift_Reg_output_3, S0=>nx14774);
   ix6812 : mux21_ni port map ( Y=>nx6811, A0=>
      booth_integrtaion_2_shift_Reg_count_3, A1=>
      booth_integrtaion_2_shift_Reg_output_3, S0=>nx14642);
   ix6802 : mux21_ni port map ( Y=>nx6801, A0=>
      booth_integrtaion_2_shift_Reg_count_3, A1=>
      booth_integrtaion_2_shift_Reg_output_2, S0=>nx14774);
   ix6792 : mux21_ni port map ( Y=>nx6791, A0=>
      booth_integrtaion_2_shift_Reg_count_2, A1=>
      booth_integrtaion_2_shift_Reg_output_2, S0=>nx14642);
   ix6782 : mux21_ni port map ( Y=>nx6781, A0=>
      booth_integrtaion_2_shift_Reg_count_2, A1=>
      booth_integrtaion_2_shift_Reg_output_1, S0=>nx14774);
   ix6772 : mux21_ni port map ( Y=>nx6771, A0=>
      booth_integrtaion_2_shift_Reg_count_1, A1=>
      booth_integrtaion_2_shift_Reg_output_1, S0=>nx14642);
   ix6762 : mux21_ni port map ( Y=>nx6761, A0=>
      booth_integrtaion_2_shift_Reg_count_1, A1=>nx14328, S0=>nx14776);
   ix7009 : and02 port map ( Y=>nx7008, A0=>nx12670, A1=>
      booth_integration_output_2_0);
   ix12673 : or03 port map ( Y=>nx12672, A0=>nx12549, A1=>
      booth_integrtaion_2_shift_reg_output_0, A2=>nx14850);
   ix7092 : mux21_ni port map ( Y=>nx7091, A0=>
      booth_integrtaion_2_booth_output_16, A1=>nx7538, S0=>nx14776);
   ix7539 : nor02ii port map ( Y=>nx7538, A0=>nx12680, A1=>nx14782);
   ix7015 : nor02ii port map ( Y=>nx7014, A0=>nx12665, A1=>
      booth_integrtaion_2_booth_output_16);
   ix7533 : xor2 port map ( Y=>nx2970, A0=>nx12686, A1=>nx12962);
   ix7521 : xor2 port map ( Y=>nx2971, A0=>nx12700, A1=>nx14554);
   ix7062 : mux21_ni port map ( Y=>nx7061, A0=>
      booth_integrtaion_2_booth_output_19, A1=>nx7502, S0=>nx14776);
   ix7503 : nor02ii port map ( Y=>nx7502, A0=>nx12718, A1=>nx14782);
   ix12732 : nor02_2x port map ( Y=>nx7004, A0=>nx12670, A1=>
      booth_integration_output_2_0);
   ix12735 : xor2 port map ( Y=>nx12734, A0=>nx12738, A1=>nx7110);
   ix7042 : mux21_ni port map ( Y=>nx7041, A0=>
      booth_integrtaion_2_booth_output_21, A1=>nx7478, S0=>nx14776);
   ix7479 : nor02ii port map ( Y=>nx7478, A0=>nx12758, A1=>nx14782);
   ix12771 : xor2 port map ( Y=>nx12770, A0=>nx12774, A1=>nx7158);
   ix7022 : mux21_ni port map ( Y=>nx7021, A0=>
      booth_integrtaion_2_booth_output_23, A1=>nx7454, S0=>nx14776);
   ix7455 : nor02ii port map ( Y=>nx7454, A0=>nx12794, A1=>nx14782);
   ix12807 : xor2 port map ( Y=>nx12806, A0=>nx12810, A1=>nx7206);
   ix7002 : mux21_ni port map ( Y=>nx7001, A0=>
      booth_integrtaion_2_booth_output_25, A1=>nx7430, S0=>nx14776);
   ix7431 : nor02ii port map ( Y=>nx7430, A0=>nx12830, A1=>nx14784);
   ix12843 : xor2 port map ( Y=>nx12842, A0=>nx12846, A1=>nx7254);
   ix6982 : mux21_ni port map ( Y=>nx6981, A0=>
      booth_integrtaion_2_booth_output_27, A1=>nx7406, S0=>nx14776);
   ix7407 : nor02ii port map ( Y=>nx7406, A0=>nx12866, A1=>nx14784);
   ix12879 : xor2 port map ( Y=>nx12878, A0=>nx12882, A1=>nx7302);
   ix6962 : mux21_ni port map ( Y=>nx6961, A0=>
      booth_integrtaion_2_booth_output_29, A1=>nx7382, S0=>nx14546);
   ix7383 : nor02ii port map ( Y=>nx7382, A0=>nx12902, A1=>nx14784);
   ix12915 : xor2 port map ( Y=>nx12914, A0=>nx12922, A1=>nx7350);
   ix6952 : mux21_ni port map ( Y=>nx6951, A0=>
      booth_integrtaion_2_booth_output_31, A1=>nx7370, S0=>nx14546);
   ix7371 : nor02ii port map ( Y=>nx7370, A0=>nx12919, A1=>nx14784);
   ix7365 : xor2 port map ( Y=>nx7364, A0=>nx12922, A1=>nx12934);
   ix7551 : nor02ii port map ( Y=>nx7550, A0=>nx7014, A1=>nx14784);
   ix12992 : xor2 port map ( Y=>nx12991, A0=>nx12980, A1=>adderInput_2(2));
   ix13004 : xor2 port map ( Y=>nx13003, A0=>nx12978, A1=>adderInput_2(4));
   ix13016 : xor2 port map ( Y=>nx13015, A0=>nx12976, A1=>adderInput_2(6));
   ix13028 : xor2 port map ( Y=>nx13027, A0=>nx12974, A1=>adderInput_2(8));
   ix13040 : xor2 port map ( Y=>nx13039, A0=>nx12972, A1=>adderInput_2(10));
   ix13052 : xor2 port map ( Y=>nx13051, A0=>nx12970, A1=>adderInput_2(12));
   ix13064 : xor2 port map ( Y=>nx13063, A0=>nx12968, A1=>adderInput_2(14));
   ix13070 : xor2 port map ( Y=>nx13069, A0=>nx12966, A1=>adderInput_2(15));
   ix8879 : xor2 port map ( Y=>label_1(0), A0=>adderInput_1(0), A1=>
      booth_integration_output_1_0);
   ix7782 : mux21_ni port map ( Y=>nx7781, A0=>booth_integration_output_1_0, 
      A1=>nx8722, S0=>nx14570);
   ix8723 : mux21_ni port map ( Y=>nx8722, A0=>neuron(0), A1=>
      booth_integration_output_1_1, S0=>nx14794);
   ix7772 : mux21_ni port map ( Y=>nx7771, A0=>booth_integration_output_1_1, 
      A1=>nx8710, S0=>nx14570);
   ix8711 : mux21_ni port map ( Y=>nx8710, A0=>neuron(1), A1=>
      booth_integration_output_1_2, S0=>nx14794);
   ix7762 : mux21_ni port map ( Y=>nx7761, A0=>booth_integration_output_1_2, 
      A1=>nx8698, S0=>nx14570);
   ix8699 : mux21_ni port map ( Y=>nx8698, A0=>neuron(2), A1=>
      booth_integration_output_1_3, S0=>nx14794);
   ix7752 : mux21_ni port map ( Y=>nx7751, A0=>booth_integration_output_1_3, 
      A1=>nx8686, S0=>nx14570);
   ix8687 : mux21_ni port map ( Y=>nx8686, A0=>neuron(3), A1=>
      booth_integration_output_1_4, S0=>nx14794);
   ix7742 : mux21_ni port map ( Y=>nx7741, A0=>booth_integration_output_1_4, 
      A1=>nx8674, S0=>nx14570);
   ix8675 : mux21_ni port map ( Y=>nx8674, A0=>neuron(4), A1=>
      booth_integration_output_1_5, S0=>nx14794);
   ix7732 : mux21_ni port map ( Y=>nx7731, A0=>booth_integration_output_1_5, 
      A1=>nx8662, S0=>nx14570);
   ix8663 : mux21_ni port map ( Y=>nx8662, A0=>neuron(5), A1=>
      booth_integration_output_1_6, S0=>nx14796);
   ix7722 : mux21_ni port map ( Y=>nx7721, A0=>booth_integration_output_1_6, 
      A1=>nx8650, S0=>nx14570);
   ix8651 : mux21_ni port map ( Y=>nx8650, A0=>neuron(6), A1=>
      booth_integration_output_1_7, S0=>nx14796);
   ix7712 : mux21_ni port map ( Y=>nx7711, A0=>booth_integration_output_1_7, 
      A1=>nx8638, S0=>nx14786);
   ix8639 : mux21_ni port map ( Y=>nx8638, A0=>neuron(7), A1=>
      booth_integration_output_1_8, S0=>nx14796);
   ix7702 : mux21_ni port map ( Y=>nx7701, A0=>booth_integration_output_1_8, 
      A1=>nx8626, S0=>nx14786);
   ix8627 : mux21_ni port map ( Y=>nx8626, A0=>neuron(8), A1=>
      booth_integration_output_1_9, S0=>nx14796);
   ix7692 : mux21_ni port map ( Y=>nx7691, A0=>booth_integration_output_1_9, 
      A1=>nx8614, S0=>nx14786);
   ix8615 : mux21_ni port map ( Y=>nx8614, A0=>neuron(9), A1=>
      booth_integration_output_1_10, S0=>nx14796);
   ix7682 : mux21_ni port map ( Y=>nx7681, A0=>booth_integration_output_1_10, 
      A1=>nx8602, S0=>nx14788);
   ix8603 : mux21_ni port map ( Y=>nx8602, A0=>neuron(10), A1=>
      booth_integration_output_1_11, S0=>nx14796);
   ix7672 : mux21_ni port map ( Y=>nx7671, A0=>booth_integration_output_1_11, 
      A1=>nx8590, S0=>nx14788);
   ix8591 : mux21_ni port map ( Y=>nx8590, A0=>neuron(11), A1=>
      booth_integration_output_1_12, S0=>nx14796);
   ix7662 : mux21_ni port map ( Y=>nx7661, A0=>booth_integration_output_1_12, 
      A1=>nx8578, S0=>nx14788);
   ix8579 : mux21_ni port map ( Y=>nx8578, A0=>neuron(12), A1=>
      booth_integration_output_1_13, S0=>nx14798);
   ix7652 : mux21_ni port map ( Y=>nx7651, A0=>booth_integration_output_1_13, 
      A1=>nx8566, S0=>nx14788);
   ix8567 : mux21_ni port map ( Y=>nx8566, A0=>neuron(13), A1=>
      booth_integration_output_1_14, S0=>nx14798);
   ix7642 : mux21_ni port map ( Y=>nx7641, A0=>booth_integration_output_1_14, 
      A1=>nx8554, S0=>nx14788);
   ix8555 : mux21_ni port map ( Y=>nx8554, A0=>neuron(14), A1=>
      booth_integration_output_1_15, S0=>nx14798);
   ix7632 : mux21 port map ( Y=>nx7631, A0=>nx13489, A1=>nx13120, S0=>
      nx14788);
   ix7282 : mux21_ni port map ( Y=>nx7281, A0=>
      booth_integrtaion_1_shift_Reg_count_0, A1=>nx14350, S0=>nx14644);
   ix7268 : and02 port map ( Y=>nx7267, A0=>nx14854, A1=>
      booth_integrtaion_1_shift_Reg_count_0);
   ix7462 : mux21_ni port map ( Y=>nx7461, A0=>
      booth_integrtaion_1_shift_Reg_count_9, A1=>nx14336, S0=>nx14644);
   ix7452 : mux21_ni port map ( Y=>nx7451, A0=>
      booth_integrtaion_1_shift_Reg_count_9, A1=>
      booth_integrtaion_1_shift_Reg_output_8, S0=>nx14788);
   ix7442 : mux21_ni port map ( Y=>nx7441, A0=>
      booth_integrtaion_1_shift_Reg_count_8, A1=>
      booth_integrtaion_1_shift_Reg_output_8, S0=>nx14644);
   ix7432 : mux21_ni port map ( Y=>nx7431, A0=>
      booth_integrtaion_1_shift_Reg_count_8, A1=>
      booth_integrtaion_1_shift_Reg_output_7, S0=>nx14790);
   ix7422 : mux21_ni port map ( Y=>nx7421, A0=>
      booth_integrtaion_1_shift_Reg_count_7, A1=>
      booth_integrtaion_1_shift_Reg_output_7, S0=>nx14644);
   ix7412 : mux21_ni port map ( Y=>nx7411, A0=>
      booth_integrtaion_1_shift_Reg_count_7, A1=>
      booth_integrtaion_1_shift_Reg_output_6, S0=>nx14790);
   ix7402 : mux21_ni port map ( Y=>nx7401, A0=>
      booth_integrtaion_1_shift_Reg_count_6, A1=>
      booth_integrtaion_1_shift_Reg_output_6, S0=>nx14644);
   ix7392 : mux21_ni port map ( Y=>nx7391, A0=>
      booth_integrtaion_1_shift_Reg_count_6, A1=>
      booth_integrtaion_1_shift_Reg_output_5, S0=>nx14790);
   ix7382 : mux21_ni port map ( Y=>nx7381, A0=>
      booth_integrtaion_1_shift_Reg_count_5, A1=>
      booth_integrtaion_1_shift_Reg_output_5, S0=>nx14644);
   ix7372 : mux21_ni port map ( Y=>nx7371, A0=>
      booth_integrtaion_1_shift_Reg_count_5, A1=>
      booth_integrtaion_1_shift_Reg_output_4, S0=>nx14790);
   ix7362 : mux21_ni port map ( Y=>nx7361, A0=>
      booth_integrtaion_1_shift_Reg_count_4, A1=>
      booth_integrtaion_1_shift_Reg_output_4, S0=>nx14646);
   ix7352 : mux21_ni port map ( Y=>nx7351, A0=>
      booth_integrtaion_1_shift_Reg_count_4, A1=>
      booth_integrtaion_1_shift_Reg_output_3, S0=>nx14790);
   ix7342 : mux21_ni port map ( Y=>nx7341, A0=>
      booth_integrtaion_1_shift_Reg_count_3, A1=>
      booth_integrtaion_1_shift_Reg_output_3, S0=>nx14646);
   ix7332 : mux21_ni port map ( Y=>nx7331, A0=>
      booth_integrtaion_1_shift_Reg_count_3, A1=>
      booth_integrtaion_1_shift_Reg_output_2, S0=>nx14790);
   ix7322 : mux21_ni port map ( Y=>nx7321, A0=>
      booth_integrtaion_1_shift_Reg_count_2, A1=>
      booth_integrtaion_1_shift_Reg_output_2, S0=>nx14646);
   ix7312 : mux21_ni port map ( Y=>nx7311, A0=>
      booth_integrtaion_1_shift_Reg_count_2, A1=>
      booth_integrtaion_1_shift_Reg_output_1, S0=>nx14790);
   ix7302 : mux21_ni port map ( Y=>nx7301, A0=>
      booth_integrtaion_1_shift_Reg_count_1, A1=>
      booth_integrtaion_1_shift_Reg_output_1, S0=>nx14646);
   ix7292 : mux21_ni port map ( Y=>nx7291, A0=>
      booth_integrtaion_1_shift_Reg_count_1, A1=>nx14350, S0=>nx14792);
   ix7995 : and02 port map ( Y=>nx7994, A0=>nx13193, A1=>
      booth_integration_output_1_0);
   ix13196 : or03 port map ( Y=>nx13195, A0=>nx13072, A1=>
      booth_integrtaion_1_shift_reg_output_0, A2=>nx14854);
   ix7622 : mux21_ni port map ( Y=>nx7621, A0=>
      booth_integrtaion_1_booth_output_16, A1=>nx8524, S0=>nx14792);
   ix8525 : nor02ii port map ( Y=>nx8524, A0=>nx13203, A1=>nx14798);
   ix8001 : nor02ii port map ( Y=>nx8000, A0=>nx13188, A1=>
      booth_integrtaion_1_booth_output_16);
   ix8519 : xor2 port map ( Y=>nx2985, A0=>nx13209, A1=>nx13485);
   ix8507 : xor2 port map ( Y=>nx2986, A0=>nx13223, A1=>nx14576);
   ix7592 : mux21_ni port map ( Y=>nx7591, A0=>
      booth_integrtaion_1_booth_output_19, A1=>nx8488, S0=>nx14792);
   ix8489 : nor02ii port map ( Y=>nx8488, A0=>nx13241, A1=>nx14798);
   ix13255 : nor02_2x port map ( Y=>nx7990, A0=>nx13193, A1=>
      booth_integration_output_1_0);
   ix13258 : xor2 port map ( Y=>nx13257, A0=>nx13261, A1=>nx8096);
   ix7572 : mux21_ni port map ( Y=>nx7571, A0=>
      booth_integrtaion_1_booth_output_21, A1=>nx8464, S0=>nx14792);
   ix8465 : nor02ii port map ( Y=>nx8464, A0=>nx13281, A1=>nx14798);
   ix13294 : xor2 port map ( Y=>nx13293, A0=>nx13297, A1=>nx8144);
   ix7552 : mux21_ni port map ( Y=>nx7551, A0=>
      booth_integrtaion_1_booth_output_23, A1=>nx8440, S0=>nx14792);
   ix8441 : nor02ii port map ( Y=>nx8440, A0=>nx13317, A1=>nx14798);
   ix13330 : xor2 port map ( Y=>nx13329, A0=>nx13333, A1=>nx8192);
   ix7532 : mux21_ni port map ( Y=>nx7531, A0=>
      booth_integrtaion_1_booth_output_25, A1=>nx8416, S0=>nx14792);
   ix8417 : nor02ii port map ( Y=>nx8416, A0=>nx13353, A1=>nx14800);
   ix13366 : xor2 port map ( Y=>nx13365, A0=>nx13369, A1=>nx8240);
   ix7512 : mux21_ni port map ( Y=>nx7511, A0=>
      booth_integrtaion_1_booth_output_27, A1=>nx8392, S0=>nx14792);
   ix8393 : nor02ii port map ( Y=>nx8392, A0=>nx13389, A1=>nx14800);
   ix13402 : xor2 port map ( Y=>nx13401, A0=>nx13405, A1=>nx8288);
   ix7492 : mux21_ni port map ( Y=>nx7491, A0=>
      booth_integrtaion_1_booth_output_29, A1=>nx8368, S0=>nx14568);
   ix8369 : nor02ii port map ( Y=>nx8368, A0=>nx13425, A1=>nx14800);
   ix13438 : xor2 port map ( Y=>nx13437, A0=>nx13445, A1=>nx8336);
   ix7482 : mux21_ni port map ( Y=>nx7481, A0=>
      booth_integrtaion_1_booth_output_31, A1=>nx8356, S0=>nx14568);
   ix8357 : nor02ii port map ( Y=>nx8356, A0=>nx13442, A1=>nx14800);
   ix8351 : xor2 port map ( Y=>nx8350, A0=>nx13445, A1=>nx13457);
   ix8537 : nor02ii port map ( Y=>nx8536, A0=>nx8000, A1=>nx14800);
   ix13515 : xor2 port map ( Y=>nx13514, A0=>nx13503, A1=>adderInput_1(2));
   ix13527 : xor2 port map ( Y=>nx13526, A0=>nx13501, A1=>adderInput_1(4));
   ix13539 : xor2 port map ( Y=>nx13538, A0=>nx13499, A1=>adderInput_1(6));
   ix13551 : xor2 port map ( Y=>nx13550, A0=>nx13497, A1=>adderInput_1(8));
   ix13563 : xor2 port map ( Y=>nx13562, A0=>nx13495, A1=>adderInput_1(10));
   ix13575 : xor2 port map ( Y=>nx13574, A0=>nx13493, A1=>adderInput_1(12));
   ix13587 : xor2 port map ( Y=>nx13586, A0=>nx13491, A1=>adderInput_1(14));
   ix13593 : xor2 port map ( Y=>nx13592, A0=>nx13489, A1=>adderInput_1(15));
   ix9865 : xor2 port map ( Y=>label_0(0), A0=>adderInput_0(0), A1=>
      booth_integration_output_0_0);
   ix8312 : mux21_ni port map ( Y=>nx8311, A0=>booth_integration_output_0_0, 
      A1=>nx9708, S0=>nx14592);
   ix9709 : mux21_ni port map ( Y=>nx9708, A0=>neuron(0), A1=>
      booth_integration_output_0_1, S0=>nx14810);
   ix8302 : mux21_ni port map ( Y=>nx8301, A0=>booth_integration_output_0_1, 
      A1=>nx9696, S0=>nx14592);
   ix9697 : mux21_ni port map ( Y=>nx9696, A0=>neuron(1), A1=>
      booth_integration_output_0_2, S0=>nx14810);
   ix8292 : mux21_ni port map ( Y=>nx8291, A0=>booth_integration_output_0_2, 
      A1=>nx9684, S0=>nx14592);
   ix9685 : mux21_ni port map ( Y=>nx9684, A0=>neuron(2), A1=>
      booth_integration_output_0_3, S0=>nx14810);
   ix8282 : mux21_ni port map ( Y=>nx8281, A0=>booth_integration_output_0_3, 
      A1=>nx9672, S0=>nx14592);
   ix9673 : mux21_ni port map ( Y=>nx9672, A0=>neuron(3), A1=>
      booth_integration_output_0_4, S0=>nx14810);
   ix8272 : mux21_ni port map ( Y=>nx8271, A0=>booth_integration_output_0_4, 
      A1=>nx9660, S0=>nx14592);
   ix9661 : mux21_ni port map ( Y=>nx9660, A0=>neuron(4), A1=>
      booth_integration_output_0_5, S0=>nx14810);
   ix8262 : mux21_ni port map ( Y=>nx8261, A0=>booth_integration_output_0_5, 
      A1=>nx9648, S0=>nx14592);
   ix9649 : mux21_ni port map ( Y=>nx9648, A0=>neuron(5), A1=>
      booth_integration_output_0_6, S0=>nx14812);
   ix8252 : mux21_ni port map ( Y=>nx8251, A0=>booth_integration_output_0_6, 
      A1=>nx9636, S0=>nx14592);
   ix9637 : mux21_ni port map ( Y=>nx9636, A0=>neuron(6), A1=>
      booth_integration_output_0_7, S0=>nx14812);
   ix8242 : mux21_ni port map ( Y=>nx8241, A0=>booth_integration_output_0_7, 
      A1=>nx9624, S0=>nx14802);
   ix9625 : mux21_ni port map ( Y=>nx9624, A0=>neuron(7), A1=>
      booth_integration_output_0_8, S0=>nx14812);
   ix8232 : mux21_ni port map ( Y=>nx8231, A0=>booth_integration_output_0_8, 
      A1=>nx9612, S0=>nx14802);
   ix9613 : mux21_ni port map ( Y=>nx9612, A0=>neuron(8), A1=>
      booth_integration_output_0_9, S0=>nx14812);
   ix8222 : mux21_ni port map ( Y=>nx8221, A0=>booth_integration_output_0_9, 
      A1=>nx9600, S0=>nx14802);
   ix9601 : mux21_ni port map ( Y=>nx9600, A0=>neuron(9), A1=>
      booth_integration_output_0_10, S0=>nx14812);
   ix8212 : mux21_ni port map ( Y=>nx8211, A0=>booth_integration_output_0_10, 
      A1=>nx9588, S0=>nx14804);
   ix9589 : mux21_ni port map ( Y=>nx9588, A0=>neuron(10), A1=>
      booth_integration_output_0_11, S0=>nx14812);
   ix8202 : mux21_ni port map ( Y=>nx8201, A0=>booth_integration_output_0_11, 
      A1=>nx9576, S0=>nx14804);
   ix9577 : mux21_ni port map ( Y=>nx9576, A0=>neuron(11), A1=>
      booth_integration_output_0_12, S0=>nx14812);
   ix8192 : mux21_ni port map ( Y=>nx8191, A0=>booth_integration_output_0_12, 
      A1=>nx9564, S0=>nx14804);
   ix9565 : mux21_ni port map ( Y=>nx9564, A0=>neuron(12), A1=>
      booth_integration_output_0_13, S0=>nx14814);
   ix8182 : mux21_ni port map ( Y=>nx8181, A0=>booth_integration_output_0_13, 
      A1=>nx9552, S0=>nx14804);
   ix9553 : mux21_ni port map ( Y=>nx9552, A0=>neuron(13), A1=>
      booth_integration_output_0_14, S0=>nx14814);
   ix8172 : mux21_ni port map ( Y=>nx8171, A0=>booth_integration_output_0_14, 
      A1=>nx9540, S0=>nx14804);
   ix9541 : mux21_ni port map ( Y=>nx9540, A0=>neuron(14), A1=>
      booth_integration_output_0_15, S0=>nx14814);
   ix8162 : mux21 port map ( Y=>nx8161, A0=>nx14012, A1=>nx13643, S0=>
      nx14804);
   ix7812 : mux21_ni port map ( Y=>nx7811, A0=>
      booth_integrtaion_0_shift_Reg_count_0, A1=>nx14372, S0=>nx14648);
   ix7798 : and02 port map ( Y=>nx7797, A0=>nx14858, A1=>
      booth_integrtaion_0_shift_Reg_count_0);
   ix7992 : mux21_ni port map ( Y=>nx7991, A0=>
      booth_integrtaion_0_shift_Reg_count_9, A1=>nx14358, S0=>nx14648);
   ix7982 : mux21_ni port map ( Y=>nx7981, A0=>
      booth_integrtaion_0_shift_Reg_count_9, A1=>
      booth_integrtaion_0_shift_Reg_output_8, S0=>nx14804);
   ix7972 : mux21_ni port map ( Y=>nx7971, A0=>
      booth_integrtaion_0_shift_Reg_count_8, A1=>
      booth_integrtaion_0_shift_Reg_output_8, S0=>nx14648);
   ix7962 : mux21_ni port map ( Y=>nx7961, A0=>
      booth_integrtaion_0_shift_Reg_count_8, A1=>
      booth_integrtaion_0_shift_Reg_output_7, S0=>nx14806);
   ix7952 : mux21_ni port map ( Y=>nx7951, A0=>
      booth_integrtaion_0_shift_Reg_count_7, A1=>
      booth_integrtaion_0_shift_Reg_output_7, S0=>nx14648);
   ix7942 : mux21_ni port map ( Y=>nx7941, A0=>
      booth_integrtaion_0_shift_Reg_count_7, A1=>
      booth_integrtaion_0_shift_Reg_output_6, S0=>nx14806);
   ix7932 : mux21_ni port map ( Y=>nx7931, A0=>
      booth_integrtaion_0_shift_Reg_count_6, A1=>
      booth_integrtaion_0_shift_Reg_output_6, S0=>nx14648);
   ix7922 : mux21_ni port map ( Y=>nx7921, A0=>
      booth_integrtaion_0_shift_Reg_count_6, A1=>
      booth_integrtaion_0_shift_Reg_output_5, S0=>nx14806);
   ix7912 : mux21_ni port map ( Y=>nx7911, A0=>
      booth_integrtaion_0_shift_Reg_count_5, A1=>
      booth_integrtaion_0_shift_Reg_output_5, S0=>nx14648);
   ix7902 : mux21_ni port map ( Y=>nx7901, A0=>
      booth_integrtaion_0_shift_Reg_count_5, A1=>
      booth_integrtaion_0_shift_Reg_output_4, S0=>nx14806);
   ix7892 : mux21_ni port map ( Y=>nx7891, A0=>
      booth_integrtaion_0_shift_Reg_count_4, A1=>
      booth_integrtaion_0_shift_Reg_output_4, S0=>nx14650);
   ix7882 : mux21_ni port map ( Y=>nx7881, A0=>
      booth_integrtaion_0_shift_Reg_count_4, A1=>
      booth_integrtaion_0_shift_Reg_output_3, S0=>nx14806);
   ix7872 : mux21_ni port map ( Y=>nx7871, A0=>
      booth_integrtaion_0_shift_Reg_count_3, A1=>
      booth_integrtaion_0_shift_Reg_output_3, S0=>nx14650);
   ix7862 : mux21_ni port map ( Y=>nx7861, A0=>
      booth_integrtaion_0_shift_Reg_count_3, A1=>
      booth_integrtaion_0_shift_Reg_output_2, S0=>nx14806);
   ix7852 : mux21_ni port map ( Y=>nx7851, A0=>
      booth_integrtaion_0_shift_Reg_count_2, A1=>
      booth_integrtaion_0_shift_Reg_output_2, S0=>nx14650);
   ix7842 : mux21_ni port map ( Y=>nx7841, A0=>
      booth_integrtaion_0_shift_Reg_count_2, A1=>
      booth_integrtaion_0_shift_Reg_output_1, S0=>nx14806);
   ix7832 : mux21_ni port map ( Y=>nx7831, A0=>
      booth_integrtaion_0_shift_Reg_count_1, A1=>
      booth_integrtaion_0_shift_Reg_output_1, S0=>nx14650);
   ix7822 : mux21_ni port map ( Y=>nx7821, A0=>
      booth_integrtaion_0_shift_Reg_count_1, A1=>nx14372, S0=>nx14808);
   ix8981 : and02 port map ( Y=>nx8980, A0=>nx13716, A1=>
      booth_integration_output_0_0);
   ix13719 : or03 port map ( Y=>nx13718, A0=>nx13595, A1=>
      booth_integrtaion_0_shift_reg_output_0, A2=>nx14858);
   ix8152 : mux21_ni port map ( Y=>nx8151, A0=>
      booth_integrtaion_0_booth_output_16, A1=>nx9510, S0=>nx14808);
   ix9511 : nor02ii port map ( Y=>nx9510, A0=>nx13726, A1=>nx14814);
   ix8987 : nor02ii port map ( Y=>nx8986, A0=>nx13711, A1=>
      booth_integrtaion_0_booth_output_16);
   ix9505 : xor2 port map ( Y=>nx3000, A0=>nx13732, A1=>nx14008);
   ix9493 : xor2 port map ( Y=>nx3001, A0=>nx13746, A1=>nx14598);
   ix8122 : mux21_ni port map ( Y=>nx8121, A0=>
      booth_integrtaion_0_booth_output_19, A1=>nx9474, S0=>nx14808);
   ix9475 : nor02ii port map ( Y=>nx9474, A0=>nx13764, A1=>nx14814);
   ix13778 : nor02_2x port map ( Y=>nx8976, A0=>nx13716, A1=>
      booth_integration_output_0_0);
   ix13781 : xor2 port map ( Y=>nx13780, A0=>nx13784, A1=>nx9082);
   ix8102 : mux21_ni port map ( Y=>nx8101, A0=>
      booth_integrtaion_0_booth_output_21, A1=>nx9450, S0=>nx14808);
   ix9451 : nor02ii port map ( Y=>nx9450, A0=>nx13804, A1=>nx14814);
   ix13817 : xor2 port map ( Y=>nx13816, A0=>nx13820, A1=>nx9130);
   ix8082 : mux21_ni port map ( Y=>nx8081, A0=>
      booth_integrtaion_0_booth_output_23, A1=>nx9426, S0=>nx14808);
   ix9427 : nor02ii port map ( Y=>nx9426, A0=>nx13840, A1=>nx14814);
   ix13853 : xor2 port map ( Y=>nx13852, A0=>nx13856, A1=>nx9178);
   ix8062 : mux21_ni port map ( Y=>nx8061, A0=>
      booth_integrtaion_0_booth_output_25, A1=>nx9402, S0=>nx14808);
   ix9403 : nor02ii port map ( Y=>nx9402, A0=>nx13876, A1=>nx14816);
   ix13889 : xor2 port map ( Y=>nx13888, A0=>nx13892, A1=>nx9226);
   ix8042 : mux21_ni port map ( Y=>nx8041, A0=>
      booth_integrtaion_0_booth_output_27, A1=>nx9378, S0=>nx14808);
   ix9379 : nor02ii port map ( Y=>nx9378, A0=>nx13912, A1=>nx14816);
   ix13925 : xor2 port map ( Y=>nx13924, A0=>nx13928, A1=>nx9274);
   ix8022 : mux21_ni port map ( Y=>nx8021, A0=>
      booth_integrtaion_0_booth_output_29, A1=>nx9354, S0=>nx14590);
   ix9355 : nor02ii port map ( Y=>nx9354, A0=>nx13948, A1=>nx14816);
   ix13961 : xor2 port map ( Y=>nx13960, A0=>nx13968, A1=>nx9322);
   ix8012 : mux21_ni port map ( Y=>nx8011, A0=>
      booth_integrtaion_0_booth_output_31, A1=>nx9342, S0=>nx14590);
   ix9343 : nor02ii port map ( Y=>nx9342, A0=>nx13965, A1=>nx14816);
   ix9337 : xor2 port map ( Y=>nx9336, A0=>nx13968, A1=>nx13980);
   ix9523 : nor02ii port map ( Y=>nx9522, A0=>nx8986, A1=>nx14816);
   ix14038 : xor2 port map ( Y=>nx14037, A0=>nx14026, A1=>adderInput_0(2));
   ix14050 : xor2 port map ( Y=>nx14049, A0=>nx14024, A1=>adderInput_0(4));
   ix14062 : xor2 port map ( Y=>nx14061, A0=>nx14022, A1=>adderInput_0(6));
   ix14074 : xor2 port map ( Y=>nx14073, A0=>nx14020, A1=>adderInput_0(8));
   ix14086 : xor2 port map ( Y=>nx14085, A0=>nx14018, A1=>adderInput_0(10));
   ix14098 : xor2 port map ( Y=>nx14097, A0=>nx14016, A1=>adderInput_0(12));
   ix14110 : xor2 port map ( Y=>nx14109, A0=>nx14014, A1=>adderInput_0(14));
   ix14116 : xor2 port map ( Y=>nx14115, A0=>nx14012, A1=>adderInput_0(15));
   ix14611 : buf02 port map ( Y=>nx14612, A=>nx8731);
   ix14613 : buf02 port map ( Y=>nx14614, A=>nx8731);
   ix14615 : buf02 port map ( Y=>nx14616, A=>nx9423);
   ix14617 : buf02 port map ( Y=>nx14618, A=>nx9423);
   ix14619 : buf02 port map ( Y=>nx14620, A=>nx10029);
   ix14621 : buf02 port map ( Y=>nx14622, A=>nx10029);
   ix14623 : buf02 port map ( Y=>nx14624, A=>nx10552);
   ix14625 : buf02 port map ( Y=>nx14626, A=>nx10552);
   ix14627 : buf02 port map ( Y=>nx14628, A=>nx11075);
   ix14629 : buf02 port map ( Y=>nx14630, A=>nx11075);
   ix14631 : buf02 port map ( Y=>nx14632, A=>nx11598);
   ix14633 : buf02 port map ( Y=>nx14634, A=>nx11598);
   ix14635 : buf02 port map ( Y=>nx14636, A=>nx12121);
   ix14637 : buf02 port map ( Y=>nx14638, A=>nx12121);
   ix14639 : buf02 port map ( Y=>nx14640, A=>nx12644);
   ix14641 : buf02 port map ( Y=>nx14642, A=>nx12644);
   ix14643 : buf02 port map ( Y=>nx14644, A=>nx13167);
   ix14645 : buf02 port map ( Y=>nx14646, A=>nx13167);
   ix14647 : buf02 port map ( Y=>nx14648, A=>nx13690);
   ix14649 : buf02 port map ( Y=>nx14650, A=>nx13690);
   ix14651 : inv02 port map ( Y=>nx14652, A=>done_EXMPLR);
   ix14653 : inv02 port map ( Y=>nx14654, A=>done_EXMPLR);
   ix14655 : inv02 port map ( Y=>nx14656, A=>done_EXMPLR);
   ix14657 : inv02 port map ( Y=>nx14658, A=>nx14822);
   ix14659 : inv02 port map ( Y=>nx14660, A=>nx14822);
   ix14661 : inv02 port map ( Y=>nx14662, A=>nx14824);
   ix14663 : inv02 port map ( Y=>nx14664, A=>nx14824);
   ix14665 : inv02 port map ( Y=>nx14666, A=>
      booth_integrtaion_9_shift_reg_output_0);
   ix14667 : inv02 port map ( Y=>nx14668, A=>
      booth_integrtaion_9_shift_reg_output_0);
   ix14669 : inv02 port map ( Y=>nx14670, A=>
      booth_integrtaion_9_shift_reg_output_0);
   ix14671 : inv02 port map ( Y=>nx14672, A=>
      booth_integrtaion_9_shift_reg_output_0);
   ix14673 : inv02 port map ( Y=>nx14674, A=>nx14826);
   ix14675 : inv02 port map ( Y=>nx14676, A=>nx14826);
   ix14677 : inv02 port map ( Y=>nx14678, A=>nx14828);
   ix14679 : inv02 port map ( Y=>nx14680, A=>nx14828);
   ix14681 : inv02 port map ( Y=>nx14682, A=>
      booth_integrtaion_8_shift_reg_output_0);
   ix14683 : inv02 port map ( Y=>nx14684, A=>
      booth_integrtaion_8_shift_reg_output_0);
   ix14685 : inv02 port map ( Y=>nx14686, A=>
      booth_integrtaion_8_shift_reg_output_0);
   ix14687 : inv02 port map ( Y=>nx14688, A=>
      booth_integrtaion_8_shift_reg_output_0);
   ix14689 : inv02 port map ( Y=>nx14690, A=>nx14830);
   ix14691 : inv02 port map ( Y=>nx14692, A=>nx14830);
   ix14693 : inv02 port map ( Y=>nx14694, A=>nx14832);
   ix14695 : inv02 port map ( Y=>nx14696, A=>nx14832);
   ix14697 : inv02 port map ( Y=>nx14698, A=>
      booth_integrtaion_7_shift_reg_output_0);
   ix14699 : inv02 port map ( Y=>nx14700, A=>
      booth_integrtaion_7_shift_reg_output_0);
   ix14701 : inv02 port map ( Y=>nx14702, A=>
      booth_integrtaion_7_shift_reg_output_0);
   ix14703 : inv02 port map ( Y=>nx14704, A=>
      booth_integrtaion_7_shift_reg_output_0);
   ix14705 : inv02 port map ( Y=>nx14706, A=>nx14834);
   ix14707 : inv02 port map ( Y=>nx14708, A=>nx14834);
   ix14709 : inv02 port map ( Y=>nx14710, A=>nx14836);
   ix14711 : inv02 port map ( Y=>nx14712, A=>nx14836);
   ix14713 : inv02 port map ( Y=>nx14714, A=>
      booth_integrtaion_6_shift_reg_output_0);
   ix14715 : inv02 port map ( Y=>nx14716, A=>
      booth_integrtaion_6_shift_reg_output_0);
   ix14717 : inv02 port map ( Y=>nx14718, A=>
      booth_integrtaion_6_shift_reg_output_0);
   ix14719 : inv02 port map ( Y=>nx14720, A=>
      booth_integrtaion_6_shift_reg_output_0);
   ix14721 : inv02 port map ( Y=>nx14722, A=>nx14838);
   ix14723 : inv02 port map ( Y=>nx14724, A=>nx14838);
   ix14725 : inv02 port map ( Y=>nx14726, A=>nx14840);
   ix14727 : inv02 port map ( Y=>nx14728, A=>nx14840);
   ix14729 : inv02 port map ( Y=>nx14730, A=>
      booth_integrtaion_5_shift_reg_output_0);
   ix14731 : inv02 port map ( Y=>nx14732, A=>
      booth_integrtaion_5_shift_reg_output_0);
   ix14733 : inv02 port map ( Y=>nx14734, A=>
      booth_integrtaion_5_shift_reg_output_0);
   ix14735 : inv02 port map ( Y=>nx14736, A=>
      booth_integrtaion_5_shift_reg_output_0);
   ix14737 : inv02 port map ( Y=>nx14738, A=>nx14842);
   ix14739 : inv02 port map ( Y=>nx14740, A=>nx14842);
   ix14741 : inv02 port map ( Y=>nx14742, A=>nx14844);
   ix14743 : inv02 port map ( Y=>nx14744, A=>nx14844);
   ix14745 : inv02 port map ( Y=>nx14746, A=>
      booth_integrtaion_4_shift_reg_output_0);
   ix14747 : inv02 port map ( Y=>nx14748, A=>
      booth_integrtaion_4_shift_reg_output_0);
   ix14749 : inv02 port map ( Y=>nx14750, A=>
      booth_integrtaion_4_shift_reg_output_0);
   ix14751 : inv02 port map ( Y=>nx14752, A=>
      booth_integrtaion_4_shift_reg_output_0);
   ix14753 : inv02 port map ( Y=>nx14754, A=>nx14846);
   ix14755 : inv02 port map ( Y=>nx14756, A=>nx14846);
   ix14757 : inv02 port map ( Y=>nx14758, A=>nx14848);
   ix14759 : inv02 port map ( Y=>nx14760, A=>nx14848);
   ix14761 : inv02 port map ( Y=>nx14762, A=>
      booth_integrtaion_3_shift_reg_output_0);
   ix14763 : inv02 port map ( Y=>nx14764, A=>
      booth_integrtaion_3_shift_reg_output_0);
   ix14765 : inv02 port map ( Y=>nx14766, A=>
      booth_integrtaion_3_shift_reg_output_0);
   ix14767 : inv02 port map ( Y=>nx14768, A=>
      booth_integrtaion_3_shift_reg_output_0);
   ix14769 : inv02 port map ( Y=>nx14770, A=>nx14850);
   ix14771 : inv02 port map ( Y=>nx14772, A=>nx14850);
   ix14773 : inv02 port map ( Y=>nx14774, A=>nx14852);
   ix14775 : inv02 port map ( Y=>nx14776, A=>nx14852);
   ix14777 : inv02 port map ( Y=>nx14778, A=>
      booth_integrtaion_2_shift_reg_output_0);
   ix14779 : inv02 port map ( Y=>nx14780, A=>
      booth_integrtaion_2_shift_reg_output_0);
   ix14781 : inv02 port map ( Y=>nx14782, A=>
      booth_integrtaion_2_shift_reg_output_0);
   ix14783 : inv02 port map ( Y=>nx14784, A=>
      booth_integrtaion_2_shift_reg_output_0);
   ix14785 : inv02 port map ( Y=>nx14786, A=>nx14854);
   ix14787 : inv02 port map ( Y=>nx14788, A=>nx14854);
   ix14789 : inv02 port map ( Y=>nx14790, A=>nx14856);
   ix14791 : inv02 port map ( Y=>nx14792, A=>nx14856);
   ix14793 : inv02 port map ( Y=>nx14794, A=>
      booth_integrtaion_1_shift_reg_output_0);
   ix14795 : inv02 port map ( Y=>nx14796, A=>
      booth_integrtaion_1_shift_reg_output_0);
   ix14797 : inv02 port map ( Y=>nx14798, A=>
      booth_integrtaion_1_shift_reg_output_0);
   ix14799 : inv02 port map ( Y=>nx14800, A=>
      booth_integrtaion_1_shift_reg_output_0);
   ix14801 : inv02 port map ( Y=>nx14802, A=>nx14858);
   ix14803 : inv02 port map ( Y=>nx14804, A=>nx14858);
   ix14805 : inv02 port map ( Y=>nx14806, A=>nx14860);
   ix14807 : inv02 port map ( Y=>nx14808, A=>nx14860);
   ix14809 : inv02 port map ( Y=>nx14810, A=>
      booth_integrtaion_0_shift_reg_output_0);
   ix14811 : inv02 port map ( Y=>nx14812, A=>
      booth_integrtaion_0_shift_reg_output_0);
   ix14813 : inv02 port map ( Y=>nx14814, A=>
      booth_integrtaion_0_shift_reg_output_0);
   ix14815 : inv02 port map ( Y=>nx14816, A=>
      booth_integrtaion_0_shift_reg_output_0);
   ix14821 : inv02 port map ( Y=>nx14822, A=>nx14388);
   ix14823 : inv02 port map ( Y=>nx14824, A=>nx14388);
   ix14825 : inv02 port map ( Y=>nx14826, A=>nx14410);
   ix14827 : inv02 port map ( Y=>nx14828, A=>nx14410);
   ix14829 : inv02 port map ( Y=>nx14830, A=>nx14432);
   ix14831 : inv02 port map ( Y=>nx14832, A=>nx14432);
   ix14833 : inv02 port map ( Y=>nx14834, A=>nx14454);
   ix14835 : inv02 port map ( Y=>nx14836, A=>nx14454);
   ix14837 : inv02 port map ( Y=>nx14838, A=>nx14476);
   ix14839 : inv02 port map ( Y=>nx14840, A=>nx14476);
   ix14841 : inv02 port map ( Y=>nx14842, A=>nx14498);
   ix14843 : inv02 port map ( Y=>nx14844, A=>nx14498);
   ix14845 : inv02 port map ( Y=>nx14846, A=>nx14520);
   ix14847 : inv02 port map ( Y=>nx14848, A=>nx14520);
   ix14849 : inv02 port map ( Y=>nx14850, A=>nx14542);
   ix14851 : inv02 port map ( Y=>nx14852, A=>nx14542);
   ix14853 : inv02 port map ( Y=>nx14854, A=>nx14564);
   ix14855 : inv02 port map ( Y=>nx14856, A=>nx14564);
   ix14857 : inv02 port map ( Y=>nx14858, A=>nx14586);
   ix14859 : inv02 port map ( Y=>nx14860, A=>nx14586);
end my_booth_adder_components ;


