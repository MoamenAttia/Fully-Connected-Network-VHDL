//
// Verilog description for cell controller, 
// Sun Apr 21 14:19:10 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module controller ( clk, clk_inv, rst, initiate, ready_signal, done, 
                    enable_mar_in, enable_mdr_in, enable_mdr_out, enable_write, 
                    mdr_data_out, label_1_output, label_2_output, label_3_output, 
                    label_4_output, label_5_output, label_6_output, 
                    label_7_output, label_8_output, label_9_output, 
                    label_10_output, state, sub_state, answer, done_comp ) ;

    input clk ;
    input clk_inv ;
    input rst ;
    inout initiate ;
    inout ready_signal ;
    inout done ;
    inout enable_mar_in ;
    inout enable_mdr_in ;
    inout enable_mdr_out ;
    inout enable_write ;
    inout [255:0]mdr_data_out ;
    inout [15:0]label_1_output ;
    inout [15:0]label_2_output ;
    inout [15:0]label_3_output ;
    inout [15:0]label_4_output ;
    inout [15:0]label_5_output ;
    inout [15:0]label_6_output ;
    inout [15:0]label_7_output ;
    inout [15:0]label_8_output ;
    inout [15:0]label_9_output ;
    inout [15:0]label_10_output ;
    inout [2:0]state ;
    inout [2:0]sub_state ;
    output [15:0]answer ;
    inout done_comp ;

    wire sel_dst_0, nx12877, num_out_2, nx4, nx12879, nx12882, nx12883, nx12885, 
         nx12887, nx20, nx26, nx38, nx56, nx64, enable_decoder_dst_booth, 
         booth_shift_Reg_adder_0_output_17, booth_shift_Reg_adder_0_output_16, 
         booth_shift_Reg_adder_0_output_15, booth_shift_Reg_adder_0_output_14, 
         booth_shift_Reg_adder_0_output_13, booth_shift_Reg_adder_0_output_12, 
         booth_shift_Reg_adder_0_output_11, booth_shift_Reg_adder_0_output_10, 
         booth_shift_Reg_adder_0_output_9, booth_shift_Reg_adder_0_output_8, 
         booth_shift_Reg_adder_0_output_7, booth_shift_Reg_adder_0_output_6, 
         booth_shift_Reg_adder_0_output_5, booth_shift_Reg_adder_0_output_4, 
         booth_shift_Reg_adder_0_output_3, booth_shift_Reg_adder_0_output_2, 
         booth_shift_Reg_adder_0_output_1, booth_shift_Reg_adder_0_output_0, 
         nx12891, nx172, nx12893, nx174, nx186, nx190, nx210, num_in_2, nx242, 
         nx258, nx266, nx278, nx12895, alu_inp1_0, address_out_0, enable_address, 
         nx300, address_in_0, nx320, nx334, nx350, nx358, num_out_0, num_in_0, 
         nx376, nx390, nx412, alu_inp1_1, address_out_1, address_in_1, nx12898, 
         nx414, nx416, num_out_1, num_in_1, nx448, alu_inp1_2, address_out_2, 
         address_in_2, nx464, nx480, nx496, nx516, num_out_3, num_in_3, nx522, 
         alu_inp1_3, address_out_3, address_in_3, nx12901, nx524, nx540, nx548, 
         num_out_4, num_in_4, alu_inp1_4, address_out_4, address_in_4, nx574, 
         nx590, nx606, num_out_5, nx630, alu_inp1_5, address_out_5, address_in_5, 
         nx12905, nx632, nx648, nx656, num_out_6, num_in_6, alu_inp1_6, 
         address_out_6, address_in_6, nx682, nx698, nx714, num_out_7, nx736, 
         alu_inp1_7, address_out_7, address_in_7, nx12907, nx738, nx754, nx12909, 
         nx830, nx846, nx868, nx878, label_4_input_15, 
         label_4_input_state_machine_15, label_4_input_0, 
         booth_booth_integrtaion_3_shift_reg_output_9, 
         booth_booth_integrtaion_3_shift_Reg_count_9, 
         booth_booth_integrtaion_3_shift_Reg_output_8, 
         booth_booth_integrtaion_3_shift_Reg_count_8, 
         booth_booth_integrtaion_3_shift_Reg_output_7, 
         booth_booth_integrtaion_3_shift_Reg_count_7, 
         booth_booth_integrtaion_3_shift_Reg_output_6, 
         booth_booth_integrtaion_3_shift_Reg_count_6, 
         booth_booth_integrtaion_3_shift_Reg_output_5, 
         booth_booth_integrtaion_3_shift_Reg_count_5, 
         booth_booth_integrtaion_3_shift_Reg_output_4, 
         booth_booth_integrtaion_3_shift_Reg_count_4, 
         booth_booth_integrtaion_3_shift_Reg_output_3, 
         booth_booth_integrtaion_3_shift_Reg_count_3, 
         booth_booth_integrtaion_3_shift_Reg_output_2, 
         booth_booth_integrtaion_3_shift_Reg_count_2, 
         booth_booth_integrtaion_3_shift_Reg_output_1, 
         booth_booth_integrtaion_3_shift_Reg_count_1, 
         booth_booth_integrtaion_3_shift_reg_output_0, 
         booth_booth_integrtaion_3_shift_Reg_count_0, 
         booth_booth_integration_output_3_1, booth_booth_integration_output_3_2, 
         booth_booth_integration_output_3_3, booth_booth_integration_output_3_4, 
         booth_booth_integration_output_3_5, booth_booth_integration_output_3_6, 
         booth_booth_integration_output_3_7, booth_booth_integration_output_3_8, 
         booth_booth_integration_output_3_9, booth_booth_integration_output_3_10, 
         booth_booth_integration_output_3_11, 
         booth_booth_integration_output_3_12, 
         booth_booth_integration_output_3_13, 
         booth_booth_integration_output_3_14, 
         booth_booth_integration_output_3_15, 
         booth_booth_integrtaion_3_booth_output_16, nx994, nx1000, 
         booth_booth_integrtaion_3_booth_output_17, nx12913, nx1008, nx1024, 
         booth_booth_integrtaion_3_booth_output_18, nx12915, nx1034, nx1038, 
         nx1052, booth_booth_integrtaion_3_booth_output_19, nx12917, nx1058, 
         nx1062, nx1072, booth_booth_integrtaion_3_booth_output_20, nx12919, 
         nx1082, nx1086, nx1100, booth_booth_integrtaion_3_booth_output_21, 
         nx12921, nx1106, nx1110, nx1120, 
         booth_booth_integrtaion_3_booth_output_22, nx12922, nx1130, nx1134, 
         nx1148, booth_booth_integrtaion_3_booth_output_23, nx12923, nx1154, 
         nx1158, nx1168, booth_booth_integrtaion_3_booth_output_24, nx12925, 
         nx1178, nx1182, nx1196, booth_booth_integrtaion_3_booth_output_25, 
         nx12927, nx1202, nx1206, nx1216, 
         booth_booth_integrtaion_3_booth_output_26, nx12929, nx1226, nx1230, 
         nx1244, booth_booth_integrtaion_3_booth_output_27, nx12930, nx1250, 
         nx1254, nx1264, booth_booth_integrtaion_3_booth_output_28, nx12931, 
         nx1274, nx1278, nx1292, booth_booth_integrtaion_3_booth_output_29, 
         nx12933, nx1298, nx1302, nx1312, 
         booth_booth_integrtaion_3_booth_output_31, nx12935, nx1322, nx1326, 
         nx1340, nx1342, nx1350, nx1356, nx1364, nx1380, nx1388, nx1404, nx1412, 
         nx1428, nx1436, nx1452, nx1460, nx1476, nx1484, nx1500, nx1508, nx1524, 
         nx1530, nx1536, nx1554, nx1566, nx1578, nx1590, nx1602, nx1614, nx1626, 
         nx1638, nx1650, nx1662, nx1674, nx1686, nx1698, nx1710, nx1722, nx1732, 
         label_4_input_state_machine_0, nx1744, label_4_input_1, 
         label_4_input_state_machine_1, nx12939, nx1766, nx1770, label_4_input_2, 
         label_4_input_state_machine_2, nx1798, nx1802, nx1820, label_4_input_3, 
         label_4_input_state_machine_3, nx12943, nx1830, nx1834, label_4_input_4, 
         label_4_input_state_machine_4, nx1862, nx1866, nx1884, label_4_input_5, 
         label_4_input_state_machine_5, nx12946, nx1894, nx1898, label_4_input_6, 
         label_4_input_state_machine_6, nx1926, nx1930, nx1948, label_4_input_7, 
         label_4_input_state_machine_7, nx12949, nx1958, nx1962, label_4_input_8, 
         label_4_input_state_machine_8, nx1990, nx1994, nx2012, label_4_input_9, 
         label_4_input_state_machine_9, nx12953, nx2022, nx2026, 
         label_4_input_10, label_4_input_state_machine_10, nx2054, nx2058, 
         nx2076, label_4_input_11, label_4_input_state_machine_11, nx12955, 
         nx2086, nx2090, label_4_input_12, label_4_input_state_machine_12, 
         nx2118, nx2122, nx2140, label_4_input_13, 
         label_4_input_state_machine_13, nx12959, nx2150, nx2154, 
         label_4_input_14, label_4_input_state_machine_14, nx2182, nx2186, 
         nx2204, nx2208, nx2212, label_3_input_15, 
         label_3_input_state_machine_15, label_3_input_0, 
         booth_booth_integrtaion_2_shift_reg_output_9, 
         booth_booth_integrtaion_2_shift_Reg_count_9, 
         booth_booth_integrtaion_2_shift_Reg_output_8, 
         booth_booth_integrtaion_2_shift_Reg_count_8, 
         booth_booth_integrtaion_2_shift_Reg_output_7, 
         booth_booth_integrtaion_2_shift_Reg_count_7, 
         booth_booth_integrtaion_2_shift_Reg_output_6, 
         booth_booth_integrtaion_2_shift_Reg_count_6, 
         booth_booth_integrtaion_2_shift_Reg_output_5, 
         booth_booth_integrtaion_2_shift_Reg_count_5, 
         booth_booth_integrtaion_2_shift_Reg_output_4, 
         booth_booth_integrtaion_2_shift_Reg_count_4, 
         booth_booth_integrtaion_2_shift_Reg_output_3, 
         booth_booth_integrtaion_2_shift_Reg_count_3, 
         booth_booth_integrtaion_2_shift_Reg_output_2, 
         booth_booth_integrtaion_2_shift_Reg_count_2, 
         booth_booth_integrtaion_2_shift_Reg_output_1, 
         booth_booth_integrtaion_2_shift_Reg_count_1, 
         booth_booth_integrtaion_2_shift_reg_output_0, 
         booth_booth_integrtaion_2_shift_Reg_count_0, 
         booth_booth_integration_output_2_1, booth_booth_integration_output_2_2, 
         booth_booth_integration_output_2_3, booth_booth_integration_output_2_4, 
         booth_booth_integration_output_2_5, booth_booth_integration_output_2_6, 
         booth_booth_integration_output_2_7, booth_booth_integration_output_2_8, 
         booth_booth_integration_output_2_9, booth_booth_integration_output_2_10, 
         booth_booth_integration_output_2_11, 
         booth_booth_integration_output_2_12, 
         booth_booth_integration_output_2_13, 
         booth_booth_integration_output_2_14, 
         booth_booth_integration_output_2_15, 
         booth_booth_integrtaion_2_booth_output_16, nx2332, nx2338, 
         booth_booth_integrtaion_2_booth_output_17, nx12965, nx2346, nx2362, 
         booth_booth_integrtaion_2_booth_output_18, nx12967, nx2372, nx2376, 
         nx2390, booth_booth_integrtaion_2_booth_output_19, nx12969, nx2396, 
         nx2400, nx2410, booth_booth_integrtaion_2_booth_output_20, nx12970, 
         nx2420, nx2424, nx2438, booth_booth_integrtaion_2_booth_output_21, 
         nx12971, nx2444, nx2448, nx2458, 
         booth_booth_integrtaion_2_booth_output_22, nx12973, nx2468, nx2472, 
         nx2486, booth_booth_integrtaion_2_booth_output_23, nx12975, nx2492, 
         nx2496, nx2506, booth_booth_integrtaion_2_booth_output_24, nx12977, 
         nx2516, nx2520, nx2534, booth_booth_integrtaion_2_booth_output_25, 
         nx12978, nx2540, nx2544, nx2554, 
         booth_booth_integrtaion_2_booth_output_26, nx12979, nx2564, nx2568, 
         nx2582, booth_booth_integrtaion_2_booth_output_27, nx12981, nx2588, 
         nx2592, nx2602, booth_booth_integrtaion_2_booth_output_28, nx12983, 
         nx2612, nx2616, nx2630, booth_booth_integrtaion_2_booth_output_29, 
         nx12985, nx2636, nx2640, nx2650, 
         booth_booth_integrtaion_2_booth_output_31, nx12987, nx2660, nx2664, 
         nx2678, nx2680, nx2688, nx2694, nx2702, nx2718, nx2726, nx2742, nx2750, 
         nx2766, nx2774, nx2790, nx2798, nx2814, nx2822, nx2838, nx2846, nx2862, 
         nx2868, nx2874, nx2892, nx2904, nx2916, nx2928, nx2940, nx2952, nx2964, 
         nx2976, nx2988, nx3000, nx3012, nx3024, nx3036, nx3048, nx3060, nx3070, 
         label_3_input_state_machine_0, nx3082, label_3_input_1, 
         label_3_input_state_machine_1, nx12991, nx3104, nx3108, label_3_input_2, 
         label_3_input_state_machine_2, nx3136, nx3140, nx3158, label_3_input_3, 
         label_3_input_state_machine_3, nx12994, nx3168, nx3172, label_3_input_4, 
         label_3_input_state_machine_4, nx3200, nx3204, nx3222, label_3_input_5, 
         label_3_input_state_machine_5, nx12997, nx3232, nx3236, label_3_input_6, 
         label_3_input_state_machine_6, nx3264, nx3268, nx3286, label_3_input_7, 
         label_3_input_state_machine_7, nx13001, nx3296, nx3300, label_3_input_8, 
         label_3_input_state_machine_8, nx3328, nx3332, nx3350, label_3_input_9, 
         label_3_input_state_machine_9, nx13003, nx3360, nx3364, 
         label_3_input_10, label_3_input_state_machine_10, nx3392, nx3396, 
         nx3414, label_3_input_11, label_3_input_state_machine_11, nx13007, 
         nx3424, nx3428, label_3_input_12, label_3_input_state_machine_12, 
         nx3456, nx3460, nx3478, label_3_input_13, 
         label_3_input_state_machine_13, nx13011, nx3488, nx3492, 
         label_3_input_14, label_3_input_state_machine_14, nx3520, nx3524, 
         nx3542, nx3546, nx3550, label_2_input_15, 
         label_2_input_state_machine_15, label_2_input_0, 
         booth_booth_integrtaion_1_shift_reg_output_9, 
         booth_booth_integrtaion_1_shift_Reg_count_9, 
         booth_booth_integrtaion_1_shift_Reg_output_8, 
         booth_booth_integrtaion_1_shift_Reg_count_8, 
         booth_booth_integrtaion_1_shift_Reg_output_7, 
         booth_booth_integrtaion_1_shift_Reg_count_7, 
         booth_booth_integrtaion_1_shift_Reg_output_6, 
         booth_booth_integrtaion_1_shift_Reg_count_6, 
         booth_booth_integrtaion_1_shift_Reg_output_5, 
         booth_booth_integrtaion_1_shift_Reg_count_5, 
         booth_booth_integrtaion_1_shift_Reg_output_4, 
         booth_booth_integrtaion_1_shift_Reg_count_4, 
         booth_booth_integrtaion_1_shift_Reg_output_3, 
         booth_booth_integrtaion_1_shift_Reg_count_3, 
         booth_booth_integrtaion_1_shift_Reg_output_2, 
         booth_booth_integrtaion_1_shift_Reg_count_2, 
         booth_booth_integrtaion_1_shift_Reg_output_1, 
         booth_booth_integrtaion_1_shift_Reg_count_1, 
         booth_booth_integrtaion_1_shift_reg_output_0, 
         booth_booth_integrtaion_1_shift_Reg_count_0, 
         booth_booth_integration_output_1_1, booth_booth_integration_output_1_2, 
         booth_booth_integration_output_1_3, booth_booth_integration_output_1_4, 
         booth_booth_integration_output_1_5, booth_booth_integration_output_1_6, 
         booth_booth_integration_output_1_7, booth_booth_integration_output_1_8, 
         booth_booth_integration_output_1_9, booth_booth_integration_output_1_10, 
         booth_booth_integration_output_1_11, 
         booth_booth_integration_output_1_12, 
         booth_booth_integration_output_1_13, 
         booth_booth_integration_output_1_14, 
         booth_booth_integration_output_1_15, 
         booth_booth_integrtaion_1_booth_output_16, nx3670, nx3676, 
         booth_booth_integrtaion_1_booth_output_17, nx13017, nx3684, nx3700, 
         booth_booth_integrtaion_1_booth_output_18, nx13018, nx3710, nx3714, 
         nx3728, booth_booth_integrtaion_1_booth_output_19, nx13019, nx3734, 
         nx3738, nx3748, booth_booth_integrtaion_1_booth_output_20, nx13021, 
         nx3758, nx3762, nx3776, booth_booth_integrtaion_1_booth_output_21, 
         nx13023, nx3782, nx3786, nx3796, 
         booth_booth_integrtaion_1_booth_output_22, nx13025, nx3806, nx3810, 
         nx3824, booth_booth_integrtaion_1_booth_output_23, nx13026, nx3830, 
         nx3834, nx3844, booth_booth_integrtaion_1_booth_output_24, nx13027, 
         nx3854, nx3858, nx3872, booth_booth_integrtaion_1_booth_output_25, 
         nx13029, nx3878, nx3882, nx3892, 
         booth_booth_integrtaion_1_booth_output_26, nx13031, nx3902, nx3906, 
         nx3920, booth_booth_integrtaion_1_booth_output_27, nx13033, nx3926, 
         nx3930, nx3940, booth_booth_integrtaion_1_booth_output_28, nx13035, 
         nx3950, nx3954, nx3968, booth_booth_integrtaion_1_booth_output_29, 
         nx13037, nx3974, nx3978, nx3988, 
         booth_booth_integrtaion_1_booth_output_31, nx13039, nx3998, nx4002, 
         nx4016, nx4018, nx4026, nx4032, nx4040, nx4056, nx4064, nx4080, nx4088, 
         nx4104, nx4112, nx4128, nx4136, nx4152, nx4160, nx4176, nx4184, nx4200, 
         nx4206, nx4212, nx4230, nx4242, nx4254, nx4266, nx4278, nx4290, nx4302, 
         nx4314, nx4326, nx4338, nx4350, nx4362, nx4374, nx4386, nx4398, nx4408, 
         label_2_input_state_machine_0, nx4420, label_2_input_1, 
         label_2_input_state_machine_1, nx13042, nx4442, nx4446, label_2_input_2, 
         label_2_input_state_machine_2, nx4474, nx4478, nx4496, label_2_input_3, 
         label_2_input_state_machine_3, nx13045, nx4506, nx4510, label_2_input_4, 
         label_2_input_state_machine_4, nx4538, nx4542, nx4560, label_2_input_5, 
         label_2_input_state_machine_5, nx13049, nx4570, nx4574, label_2_input_6, 
         label_2_input_state_machine_6, nx4602, nx4606, nx4624, label_2_input_7, 
         label_2_input_state_machine_7, nx13051, nx4634, nx4638, label_2_input_8, 
         label_2_input_state_machine_8, nx4666, nx4670, nx4688, label_2_input_9, 
         label_2_input_state_machine_9, nx13055, nx4698, nx4702, 
         label_2_input_10, label_2_input_state_machine_10, nx4730, nx4734, 
         nx4752, label_2_input_11, label_2_input_state_machine_11, nx13059, 
         nx4762, nx4766, label_2_input_12, label_2_input_state_machine_12, 
         nx4794, nx4798, nx4816, label_2_input_13, 
         label_2_input_state_machine_13, nx13063, nx4826, nx4830, 
         label_2_input_14, label_2_input_state_machine_14, nx4858, nx4862, 
         nx4880, nx4884, nx4888, label_1_input_15, 
         label_1_input_state_machine_15, label_1_input_0, 
         booth_booth_integrtaion_0_shift_reg_output_9, 
         booth_booth_integrtaion_0_shift_Reg_count_9, 
         booth_booth_integrtaion_0_shift_Reg_output_8, 
         booth_booth_integrtaion_0_shift_Reg_count_8, 
         booth_booth_integrtaion_0_shift_Reg_output_7, 
         booth_booth_integrtaion_0_shift_Reg_count_7, 
         booth_booth_integrtaion_0_shift_Reg_output_6, 
         booth_booth_integrtaion_0_shift_Reg_count_6, 
         booth_booth_integrtaion_0_shift_Reg_output_5, 
         booth_booth_integrtaion_0_shift_Reg_count_5, 
         booth_booth_integrtaion_0_shift_Reg_output_4, 
         booth_booth_integrtaion_0_shift_Reg_count_4, 
         booth_booth_integrtaion_0_shift_Reg_output_3, 
         booth_booth_integrtaion_0_shift_Reg_count_3, 
         booth_booth_integrtaion_0_shift_Reg_output_2, 
         booth_booth_integrtaion_0_shift_Reg_count_2, 
         booth_booth_integrtaion_0_shift_Reg_output_1, 
         booth_booth_integrtaion_0_shift_Reg_count_1, 
         booth_booth_integrtaion_0_shift_reg_output_0, 
         booth_booth_integrtaion_0_shift_Reg_count_0, 
         booth_booth_integration_output_0_1, booth_booth_integration_output_0_2, 
         booth_booth_integration_output_0_3, booth_booth_integration_output_0_4, 
         booth_booth_integration_output_0_5, booth_booth_integration_output_0_6, 
         booth_booth_integration_output_0_7, booth_booth_integration_output_0_8, 
         booth_booth_integration_output_0_9, booth_booth_integration_output_0_10, 
         booth_booth_integration_output_0_11, 
         booth_booth_integration_output_0_12, 
         booth_booth_integration_output_0_13, 
         booth_booth_integration_output_0_14, 
         booth_booth_integration_output_0_15, 
         booth_booth_integrtaion_0_booth_output_16, nx5008, nx5014, 
         booth_booth_integrtaion_0_booth_output_17, nx13067, nx5022, nx5038, 
         booth_booth_integrtaion_0_booth_output_18, nx13069, nx5048, nx5052, 
         nx5066, booth_booth_integrtaion_0_booth_output_19, nx13071, nx5072, 
         nx5076, nx5086, booth_booth_integrtaion_0_booth_output_20, nx13073, 
         nx5096, nx5100, nx5114, booth_booth_integrtaion_0_booth_output_21, 
         nx13074, nx5120, nx5124, nx5134, 
         booth_booth_integrtaion_0_booth_output_22, nx13075, nx5144, nx5148, 
         nx5162, booth_booth_integrtaion_0_booth_output_23, nx13077, nx5168, 
         nx5172, nx5182, booth_booth_integrtaion_0_booth_output_24, nx13079, 
         nx5192, nx5196, nx5210, booth_booth_integrtaion_0_booth_output_25, 
         nx13081, nx5216, nx5220, nx5230, 
         booth_booth_integrtaion_0_booth_output_26, nx13083, nx5240, nx5244, 
         nx5258, booth_booth_integrtaion_0_booth_output_27, nx13085, nx5264, 
         nx5268, nx5278, booth_booth_integrtaion_0_booth_output_28, nx13087, 
         nx5288, nx5292, nx5306, booth_booth_integrtaion_0_booth_output_29, 
         nx13089, nx5312, nx5316, nx5326, 
         booth_booth_integrtaion_0_booth_output_31, nx13090, nx5336, nx5340, 
         nx5354, nx5356, nx5364, nx5370, nx5378, nx5394, nx5402, nx5418, nx5426, 
         nx5442, nx5450, nx5466, nx5474, nx5490, nx5498, nx5514, nx5522, nx5538, 
         nx5544, nx5550, nx5568, nx5580, nx5592, nx5604, nx5616, nx5628, nx5640, 
         nx5652, nx5664, nx5676, nx5688, nx5700, nx5712, nx5724, nx5736, nx5746, 
         label_1_input_state_machine_0, nx5758, label_1_input_1, 
         label_1_input_state_machine_1, nx13093, nx5780, nx5784, label_1_input_2, 
         label_1_input_state_machine_2, nx5812, nx5816, nx5834, label_1_input_3, 
         label_1_input_state_machine_3, nx13097, nx5844, nx5848, label_1_input_4, 
         label_1_input_state_machine_4, nx5876, nx5880, nx5898, label_1_input_5, 
         label_1_input_state_machine_5, nx13099, nx5908, nx5912, label_1_input_6, 
         label_1_input_state_machine_6, nx5940, nx5944, nx5962, label_1_input_7, 
         label_1_input_state_machine_7, nx13103, nx5972, nx5976, label_1_input_8, 
         label_1_input_state_machine_8, nx6004, nx6008, nx6026, label_1_input_9, 
         label_1_input_state_machine_9, nx13107, nx6036, nx6040, 
         label_1_input_10, label_1_input_state_machine_10, nx6068, nx6072, 
         nx6090, label_1_input_11, label_1_input_state_machine_11, nx13111, 
         nx6100, nx6104, label_1_input_12, label_1_input_state_machine_12, 
         nx6132, nx6136, nx6154, label_1_input_13, 
         label_1_input_state_machine_13, nx13114, nx6164, nx6168, 
         label_1_input_14, label_1_input_state_machine_14, nx6196, nx6200, 
         nx6218, nx6222, nx6226, max_calc_state_2, max_calc_start, start_comp, 
         nx6244, max_calc_state_0, max_calc_state_3, max_calc_state_1, nx6300, 
         nx6342, max_calc_comparator_first_inp1_0, nx6352, max_calc_ans1_0, 
         nx6368, nx13121, nx6388, max_calc_ans6_0, max_calc_ans5_0, 
         max_calc_comparator_fifth_inp1_0, label_9_input_0, 
         booth_booth_integrtaion_8_shift_reg_output_9, 
         booth_booth_integrtaion_8_shift_Reg_count_9, 
         booth_booth_integrtaion_8_shift_Reg_output_8, 
         booth_booth_integrtaion_8_shift_Reg_count_8, 
         booth_booth_integrtaion_8_shift_Reg_output_7, 
         booth_booth_integrtaion_8_shift_Reg_count_7, 
         booth_booth_integrtaion_8_shift_Reg_output_6, 
         booth_booth_integrtaion_8_shift_Reg_count_6, 
         booth_booth_integrtaion_8_shift_Reg_output_5, 
         booth_booth_integrtaion_8_shift_Reg_count_5, 
         booth_booth_integrtaion_8_shift_Reg_output_4, 
         booth_booth_integrtaion_8_shift_Reg_count_4, 
         booth_booth_integrtaion_8_shift_Reg_output_3, 
         booth_booth_integrtaion_8_shift_Reg_count_3, 
         booth_booth_integrtaion_8_shift_Reg_output_2, 
         booth_booth_integrtaion_8_shift_Reg_count_2, 
         booth_booth_integrtaion_8_shift_Reg_output_1, 
         booth_booth_integrtaion_8_shift_Reg_count_1, 
         booth_booth_integrtaion_8_shift_reg_output_0, 
         booth_booth_integrtaion_8_shift_Reg_count_0, 
         booth_booth_integration_output_8_1, booth_booth_integration_output_8_2, 
         booth_booth_integration_output_8_3, booth_booth_integration_output_8_4, 
         booth_booth_integration_output_8_5, booth_booth_integration_output_8_6, 
         booth_booth_integration_output_8_7, booth_booth_integration_output_8_8, 
         booth_booth_integration_output_8_9, booth_booth_integration_output_8_10, 
         booth_booth_integration_output_8_11, 
         booth_booth_integration_output_8_12, 
         booth_booth_integration_output_8_13, 
         booth_booth_integration_output_8_14, 
         booth_booth_integration_output_8_15, 
         booth_booth_integrtaion_8_booth_output_16, nx6508, nx6514, 
         booth_booth_integrtaion_8_booth_output_17, nx13123, nx6522, nx6538, 
         booth_booth_integrtaion_8_booth_output_18, nx13125, nx6548, nx6552, 
         nx6566, booth_booth_integrtaion_8_booth_output_19, nx13127, nx6572, 
         nx6576, nx6586, booth_booth_integrtaion_8_booth_output_20, nx13129, 
         nx6596, nx6600, nx6614, booth_booth_integrtaion_8_booth_output_21, 
         nx13131, nx6620, nx6624, nx6634, 
         booth_booth_integrtaion_8_booth_output_22, nx13133, nx6644, nx6648, 
         nx6662, booth_booth_integrtaion_8_booth_output_23, nx13135, nx6668, 
         nx6672, nx6682, booth_booth_integrtaion_8_booth_output_24, nx13137, 
         nx6692, nx6696, nx6710, booth_booth_integrtaion_8_booth_output_25, 
         nx13138, nx6716, nx6720, nx6730, 
         booth_booth_integrtaion_8_booth_output_26, nx13139, nx6740, nx6744, 
         nx6758, booth_booth_integrtaion_8_booth_output_27, nx13141, nx6764, 
         nx6768, nx6778, booth_booth_integrtaion_8_booth_output_28, nx13143, 
         nx6788, nx6792, nx6806, booth_booth_integrtaion_8_booth_output_29, 
         nx13145, nx6812, nx6816, nx6826, 
         booth_booth_integrtaion_8_booth_output_31, nx13146, nx6836, nx6840, 
         nx6854, nx6856, nx6864, nx6870, nx6878, nx6894, nx6902, nx6918, nx6926, 
         nx6942, nx6950, nx6966, nx6974, nx6990, nx6998, nx7014, nx7022, nx7038, 
         nx7044, nx7050, nx7068, nx7080, nx7092, nx7104, nx7116, nx7128, nx7140, 
         nx7152, nx7164, nx7176, nx7188, nx7200, nx7212, nx7224, nx7236, nx7248, 
         label_9_input_state_machine_0, nx7260, label_10_input_14, 
         label_10_input_state_machine_14, label_10_input_0, 
         booth_booth_integrtaion_9_shift_reg_output_9, 
         booth_booth_integrtaion_9_shift_Reg_count_9, 
         booth_booth_integrtaion_9_shift_Reg_output_8, 
         booth_booth_integrtaion_9_shift_Reg_count_8, 
         booth_booth_integrtaion_9_shift_Reg_output_7, 
         booth_booth_integrtaion_9_shift_Reg_count_7, 
         booth_booth_integrtaion_9_shift_Reg_output_6, 
         booth_booth_integrtaion_9_shift_Reg_count_6, 
         booth_booth_integrtaion_9_shift_Reg_output_5, 
         booth_booth_integrtaion_9_shift_Reg_count_5, 
         booth_booth_integrtaion_9_shift_Reg_output_4, 
         booth_booth_integrtaion_9_shift_Reg_count_4, 
         booth_booth_integrtaion_9_shift_Reg_output_3, 
         booth_booth_integrtaion_9_shift_Reg_count_3, 
         booth_booth_integrtaion_9_shift_Reg_output_2, 
         booth_booth_integrtaion_9_shift_Reg_count_2, 
         booth_booth_integrtaion_9_shift_Reg_output_1, 
         booth_booth_integrtaion_9_shift_Reg_count_1, 
         booth_booth_integrtaion_9_shift_reg_output_0, 
         booth_booth_integrtaion_9_shift_Reg_count_0, 
         booth_booth_integration_output_9_1, booth_booth_integration_output_9_2, 
         booth_booth_integration_output_9_3, booth_booth_integration_output_9_4, 
         booth_booth_integration_output_9_5, booth_booth_integration_output_9_6, 
         booth_booth_integration_output_9_7, booth_booth_integration_output_9_8, 
         booth_booth_integration_output_9_9, booth_booth_integration_output_9_10, 
         booth_booth_integration_output_9_11, 
         booth_booth_integration_output_9_12, 
         booth_booth_integration_output_9_13, 
         booth_booth_integration_output_9_14, 
         booth_booth_integration_output_9_15, 
         booth_booth_integrtaion_9_booth_output_16, nx7388, nx7394, 
         booth_booth_integrtaion_9_booth_output_17, nx13149, nx7402, nx7418, 
         booth_booth_integrtaion_9_booth_output_18, nx13151, nx7428, nx7432, 
         nx7446, booth_booth_integrtaion_9_booth_output_19, nx13153, nx7452, 
         nx7456, nx7466, booth_booth_integrtaion_9_booth_output_20, nx13155, 
         nx7476, nx7480, nx7494, booth_booth_integrtaion_9_booth_output_21, 
         nx13157, nx7500, nx7504, nx7514, 
         booth_booth_integrtaion_9_booth_output_22, nx13159, nx7524, nx7528, 
         nx7542, booth_booth_integrtaion_9_booth_output_23, nx13161, nx7548, 
         nx7552, nx7562, booth_booth_integrtaion_9_booth_output_24, nx13162, 
         nx7572, nx7576, nx7590, booth_booth_integrtaion_9_booth_output_25, 
         nx13163, nx7596, nx7600, nx7610, 
         booth_booth_integrtaion_9_booth_output_26, nx13165, nx7620, nx7624, 
         nx7638, booth_booth_integrtaion_9_booth_output_27, nx13167, nx7644, 
         nx7648, nx7658, booth_booth_integrtaion_9_booth_output_28, nx13169, 
         nx7668, nx7672, nx7686, booth_booth_integrtaion_9_booth_output_29, 
         nx13170, nx7692, nx7696, nx7706, 
         booth_booth_integrtaion_9_booth_output_31, nx13171, nx7716, nx7720, 
         nx7734, nx7736, nx7744, nx7750, nx7758, nx7774, nx7782, nx7798, nx7806, 
         nx7822, nx7830, nx7846, nx7854, nx7870, nx7878, nx7894, nx7902, nx7918, 
         nx7924, nx7930, nx7948, nx7960, nx7972, nx7984, nx7996, nx8008, nx8020, 
         nx8032, nx8044, nx8056, nx8068, nx8080, nx8092, nx8104, nx8116, nx8126, 
         label_10_input_state_machine_0, nx8138, label_10_input_1, 
         label_10_input_state_machine_1, nx13175, nx8160, nx8164, 
         label_10_input_2, label_10_input_state_machine_2, nx8192, nx8196, 
         nx8214, label_10_input_3, label_10_input_state_machine_3, nx13179, 
         nx8224, nx8228, label_10_input_4, label_10_input_state_machine_4, 
         nx8256, nx8260, nx8278, label_10_input_5, 
         label_10_input_state_machine_5, nx13183, nx8288, nx8292, 
         label_10_input_6, label_10_input_state_machine_6, nx8320, nx8324, 
         nx8342, label_10_input_7, label_10_input_state_machine_7, nx13187, 
         nx8352, nx8356, label_10_input_8, label_10_input_state_machine_8, 
         nx8384, nx8388, nx8406, label_10_input_9, 
         label_10_input_state_machine_9, nx13191, nx8416, nx8420, 
         label_10_input_10, label_10_input_state_machine_10, nx8448, nx8452, 
         nx8470, label_10_input_11, label_10_input_state_machine_11, nx13195, 
         nx8480, nx8484, label_10_input_12, label_10_input_state_machine_12, 
         nx8512, nx8516, nx8534, label_10_input_13, 
         label_10_input_state_machine_13, nx13199, nx8544, nx8548, nx8570, 
         nx8574, max_calc_comparator_fifth_inp1_14, label_9_input_14, 
         label_9_input_state_machine_14, label_9_input_1, 
         label_9_input_state_machine_1, nx13200, nx8610, nx8614, label_9_input_2, 
         label_9_input_state_machine_2, nx8642, nx8646, nx8664, label_9_input_3, 
         label_9_input_state_machine_3, nx13202, nx8674, nx8678, label_9_input_4, 
         label_9_input_state_machine_4, nx8706, nx8710, nx8728, label_9_input_5, 
         label_9_input_state_machine_5, nx13204, nx8738, nx8742, label_9_input_6, 
         label_9_input_state_machine_6, nx8770, nx8774, nx8792, label_9_input_7, 
         label_9_input_state_machine_7, nx13207, nx8802, nx8806, label_9_input_8, 
         label_9_input_state_machine_8, nx8834, nx8838, nx8856, label_9_input_9, 
         label_9_input_state_machine_9, nx13211, nx8866, nx8870, 
         label_9_input_10, label_9_input_state_machine_10, nx8898, nx8902, 
         nx8920, label_9_input_11, label_9_input_state_machine_11, nx13213, 
         nx8930, nx8934, label_9_input_12, label_9_input_state_machine_12, 
         nx8962, nx8966, nx8984, label_9_input_13, 
         label_9_input_state_machine_13, nx13215, nx8994, nx8998, nx9020, nx9024, 
         nx9044, max_calc_comparator_fifth_inp2_13, 
         max_calc_comparator_fifth_inp1_13, max_calc_comparator_fifth_inp1_12, 
         nx9080, max_calc_comparator_fifth_inp2_11, 
         max_calc_comparator_fifth_inp1_11, max_calc_comparator_fifth_inp1_10, 
         nx9116, max_calc_comparator_fifth_inp2_9, 
         max_calc_comparator_fifth_inp1_9, max_calc_comparator_fifth_inp1_8, 
         nx9152, max_calc_comparator_fifth_inp2_7, 
         max_calc_comparator_fifth_inp1_7, max_calc_comparator_fifth_inp1_6, 
         nx9188, max_calc_comparator_fifth_inp2_5, 
         max_calc_comparator_fifth_inp1_5, max_calc_comparator_fifth_inp1_4, 
         nx9224, max_calc_comparator_fifth_inp2_3, 
         max_calc_comparator_fifth_inp1_3, max_calc_comparator_fifth_inp1_2, 
         nx9260, max_calc_comparator_fifth_inp2_1, nx9278, nx9302, nx9318, 
         nx9334, nx9350, nx9366, nx9382, nx9398, label_10_input_15, 
         label_10_input_state_machine_15, nx9420, nx9424, nx9428, 
         label_9_input_15, label_9_input_state_machine_15, nx9460, nx9464, 
         nx9468, nx9488, nx9490, nx9498, nx9508, nx9512, 
         max_calc_comparator_first_inp2_14, max_calc_ans2_14, 
         max_calc_comparator_second_inp1_14, max_calc_ans3_14, 
         max_calc_comparator_third_inp1_14, label_5_input_14, 
         label_5_input_state_machine_14, label_5_input_0, 
         booth_booth_integrtaion_4_shift_reg_output_9, 
         booth_booth_integrtaion_4_shift_Reg_count_9, 
         booth_booth_integrtaion_4_shift_Reg_output_8, 
         booth_booth_integrtaion_4_shift_Reg_count_8, 
         booth_booth_integrtaion_4_shift_Reg_output_7, 
         booth_booth_integrtaion_4_shift_Reg_count_7, 
         booth_booth_integrtaion_4_shift_Reg_output_6, 
         booth_booth_integrtaion_4_shift_Reg_count_6, 
         booth_booth_integrtaion_4_shift_Reg_output_5, 
         booth_booth_integrtaion_4_shift_Reg_count_5, 
         booth_booth_integrtaion_4_shift_Reg_output_4, 
         booth_booth_integrtaion_4_shift_Reg_count_4, 
         booth_booth_integrtaion_4_shift_Reg_output_3, 
         booth_booth_integrtaion_4_shift_Reg_count_3, 
         booth_booth_integrtaion_4_shift_Reg_output_2, 
         booth_booth_integrtaion_4_shift_Reg_count_2, 
         booth_booth_integrtaion_4_shift_Reg_output_1, 
         booth_booth_integrtaion_4_shift_Reg_count_1, 
         booth_booth_integrtaion_4_shift_reg_output_0, 
         booth_booth_integrtaion_4_shift_Reg_count_0, 
         booth_booth_integration_output_4_1, booth_booth_integration_output_4_2, 
         booth_booth_integration_output_4_3, booth_booth_integration_output_4_4, 
         booth_booth_integration_output_4_5, booth_booth_integration_output_4_6, 
         booth_booth_integration_output_4_7, booth_booth_integration_output_4_8, 
         booth_booth_integration_output_4_9, booth_booth_integration_output_4_10, 
         booth_booth_integration_output_4_11, 
         booth_booth_integration_output_4_12, 
         booth_booth_integration_output_4_13, 
         booth_booth_integration_output_4_14, 
         booth_booth_integration_output_4_15, 
         booth_booth_integrtaion_4_booth_output_16, nx9646, nx9652, 
         booth_booth_integrtaion_4_booth_output_17, nx13217, nx9660, nx9676, 
         booth_booth_integrtaion_4_booth_output_18, nx13219, nx9686, nx9690, 
         nx9704, booth_booth_integrtaion_4_booth_output_19, nx13221, nx9710, 
         nx9714, nx9724, booth_booth_integrtaion_4_booth_output_20, nx13223, 
         nx9734, nx9738, nx9752, booth_booth_integrtaion_4_booth_output_21, 
         nx13224, nx9758, nx9762, nx9772, 
         booth_booth_integrtaion_4_booth_output_22, nx13225, nx9782, nx9786, 
         nx9800, booth_booth_integrtaion_4_booth_output_23, nx13226, nx9806, 
         nx9810, nx9820, booth_booth_integrtaion_4_booth_output_24, nx13227, 
         nx9830, nx9834, nx9848, booth_booth_integrtaion_4_booth_output_25, 
         nx13228, nx9854, nx9858, nx9868, 
         booth_booth_integrtaion_4_booth_output_26, nx13229, nx9878, nx9882, 
         nx9896, booth_booth_integrtaion_4_booth_output_27, nx13231, nx9902, 
         nx9906, nx9916, booth_booth_integrtaion_4_booth_output_28, nx13233, 
         nx9926, nx9930, nx9944, booth_booth_integrtaion_4_booth_output_29, 
         nx13235, nx9950, nx9954, nx9964, 
         booth_booth_integrtaion_4_booth_output_31, nx13236, nx9974, nx9978, 
         nx9992, nx9994, nx10002, nx10008, nx10016, nx10032, nx10040, nx10056, 
         nx10064, nx10080, nx10088, nx10104, nx10112, nx10128, nx10136, nx10152, 
         nx10160, nx10176, nx10182, nx10188, nx10206, nx10218, nx10230, nx10242, 
         nx10254, nx10266, nx10278, nx10290, nx10302, nx10314, nx10326, nx10338, 
         nx10350, nx10362, nx10374, nx10384, label_5_input_state_machine_0, 
         nx10396, label_5_input_1, label_5_input_state_machine_1, nx13238, 
         nx10418, nx10422, label_5_input_2, label_5_input_state_machine_2, 
         nx10450, nx10454, nx10472, label_5_input_3, 
         label_5_input_state_machine_3, nx13240, nx10482, nx10486, 
         label_5_input_4, label_5_input_state_machine_4, nx10514, nx10518, 
         nx10536, label_5_input_5, label_5_input_state_machine_5, nx13243, 
         nx10546, nx10550, label_5_input_6, label_5_input_state_machine_6, 
         nx10578, nx10582, nx10600, label_5_input_7, 
         label_5_input_state_machine_7, nx13247, nx10610, nx10614, 
         label_5_input_8, label_5_input_state_machine_8, nx10642, nx10646, 
         nx10664, label_5_input_9, label_5_input_state_machine_9, nx13249, 
         nx10674, nx10678, label_5_input_10, label_5_input_state_machine_10, 
         nx10706, nx10710, nx10728, label_5_input_11, 
         label_5_input_state_machine_11, nx13251, nx10738, nx10742, 
         label_5_input_12, label_5_input_state_machine_12, nx10770, nx10774, 
         nx10792, label_5_input_13, label_5_input_state_machine_13, nx13253, 
         nx10802, nx10806, nx10828, nx10832, label_6_input_14, 
         label_6_input_state_machine_14, label_6_input_0, 
         booth_booth_integrtaion_5_shift_reg_output_9, 
         booth_booth_integrtaion_5_shift_Reg_count_9, 
         booth_booth_integrtaion_5_shift_Reg_output_8, 
         booth_booth_integrtaion_5_shift_Reg_count_8, 
         booth_booth_integrtaion_5_shift_Reg_output_7, 
         booth_booth_integrtaion_5_shift_Reg_count_7, 
         booth_booth_integrtaion_5_shift_Reg_output_6, 
         booth_booth_integrtaion_5_shift_Reg_count_6, 
         booth_booth_integrtaion_5_shift_Reg_output_5, 
         booth_booth_integrtaion_5_shift_Reg_count_5, 
         booth_booth_integrtaion_5_shift_Reg_output_4, 
         booth_booth_integrtaion_5_shift_Reg_count_4, 
         booth_booth_integrtaion_5_shift_Reg_output_3, 
         booth_booth_integrtaion_5_shift_Reg_count_3, 
         booth_booth_integrtaion_5_shift_Reg_output_2, 
         booth_booth_integrtaion_5_shift_Reg_count_2, 
         booth_booth_integrtaion_5_shift_Reg_output_1, 
         booth_booth_integrtaion_5_shift_Reg_count_1, 
         booth_booth_integrtaion_5_shift_reg_output_0, 
         booth_booth_integrtaion_5_shift_Reg_count_0, 
         booth_booth_integration_output_5_1, booth_booth_integration_output_5_2, 
         booth_booth_integration_output_5_3, booth_booth_integration_output_5_4, 
         booth_booth_integration_output_5_5, booth_booth_integration_output_5_6, 
         booth_booth_integration_output_5_7, booth_booth_integration_output_5_8, 
         booth_booth_integration_output_5_9, booth_booth_integration_output_5_10, 
         booth_booth_integration_output_5_11, 
         booth_booth_integration_output_5_12, 
         booth_booth_integration_output_5_13, 
         booth_booth_integration_output_5_14, 
         booth_booth_integration_output_5_15, 
         booth_booth_integrtaion_5_booth_output_16, nx10968, nx10974, 
         booth_booth_integrtaion_5_booth_output_17, nx13257, nx10982, nx10998, 
         booth_booth_integrtaion_5_booth_output_18, nx13259, nx11008, nx11012, 
         nx11026, booth_booth_integrtaion_5_booth_output_19, nx13260, nx11032, 
         nx11036, nx11046, booth_booth_integrtaion_5_booth_output_20, nx13261, 
         nx11056, nx11060, nx11074, booth_booth_integrtaion_5_booth_output_21, 
         nx13262, nx11080, nx11084, nx11094, 
         booth_booth_integrtaion_5_booth_output_22, nx13263, nx11104, nx11108, 
         nx11122, booth_booth_integrtaion_5_booth_output_23, nx13264, nx11128, 
         nx11132, nx11142, booth_booth_integrtaion_5_booth_output_24, nx13265, 
         nx11152, nx11156, nx11170, booth_booth_integrtaion_5_booth_output_25, 
         nx13267, nx11176, nx11180, nx11190, 
         booth_booth_integrtaion_5_booth_output_26, nx13269, nx11200, nx11204, 
         nx11218, booth_booth_integrtaion_5_booth_output_27, nx13271, nx11224, 
         nx11228, nx11238, booth_booth_integrtaion_5_booth_output_28, nx13272, 
         nx11248, nx11252, nx11266, booth_booth_integrtaion_5_booth_output_29, 
         nx13273, nx11272, nx11276, nx11286, 
         booth_booth_integrtaion_5_booth_output_31, nx13274, nx11296, nx11300, 
         nx11314, nx11316, nx11324, nx11330, nx11338, nx11354, nx11362, nx11378, 
         nx11386, nx11402, nx11410, nx11426, nx11434, nx11450, nx11458, nx11474, 
         nx11482, nx11498, nx11504, nx11510, nx11528, nx11540, nx11552, nx11564, 
         nx11576, nx11588, nx11600, nx11612, nx11624, nx11636, nx11648, nx11660, 
         nx11672, nx11684, nx11696, nx11706, label_6_input_state_machine_0, 
         nx11718, label_6_input_1, label_6_input_state_machine_1, nx13276, 
         nx11740, nx11744, label_6_input_2, label_6_input_state_machine_2, 
         nx11772, nx11776, nx11794, label_6_input_3, 
         label_6_input_state_machine_3, nx13279, nx11804, nx11808, 
         label_6_input_4, label_6_input_state_machine_4, nx11836, nx11840, 
         nx11858, label_6_input_5, label_6_input_state_machine_5, nx13283, 
         nx11868, nx11872, label_6_input_6, label_6_input_state_machine_6, 
         nx11900, nx11904, nx11922, label_6_input_7, 
         label_6_input_state_machine_7, nx13285, nx11932, nx11936, 
         label_6_input_8, label_6_input_state_machine_8, nx11964, nx11968, 
         nx11986, label_6_input_9, label_6_input_state_machine_9, nx13287, 
         nx11996, nx12000, label_6_input_10, label_6_input_state_machine_10, 
         nx12028, nx12032, nx12050, label_6_input_11, 
         label_6_input_state_machine_11, nx13289, nx12060, nx12064, 
         label_6_input_12, label_6_input_state_machine_12, nx12092, nx12096, 
         nx12114, label_6_input_13, label_6_input_state_machine_13, nx13293, 
         nx12124, nx12128, nx12150, nx12154, nx12176, 
         max_calc_comparator_third_inp2_13, max_calc_comparator_third_inp1_13, 
         max_calc_comparator_third_inp1_12, nx12220, 
         max_calc_comparator_third_inp2_11, max_calc_comparator_third_inp1_11, 
         max_calc_comparator_third_inp1_10, nx12264, 
         max_calc_comparator_third_inp2_9, max_calc_comparator_third_inp1_9, 
         max_calc_comparator_third_inp1_8, nx12308, 
         max_calc_comparator_third_inp2_7, max_calc_comparator_third_inp1_7, 
         max_calc_comparator_third_inp1_6, nx12352, 
         max_calc_comparator_third_inp2_5, max_calc_comparator_third_inp1_5, 
         max_calc_comparator_third_inp1_4, nx12396, 
         max_calc_comparator_third_inp2_3, max_calc_comparator_third_inp1_3, 
         max_calc_comparator_third_inp1_2, nx12440, 
         max_calc_comparator_third_inp2_1, nx12462, 
         max_calc_comparator_third_inp1_0, nx12498, nx12514, nx12530, nx12546, 
         nx12562, nx12578, nx12594, label_6_input_15, 
         label_6_input_state_machine_15, nx12616, nx12620, nx12624, 
         label_5_input_15, label_5_input_state_machine_15, nx12658, nx12662, 
         nx12666, nx12688, nx12690, nx12712, max_calc_ans4_14, 
         max_calc_comparator_fourth_inp1_14, label_7_input_14, 
         label_7_input_state_machine_14, label_7_input_0, 
         booth_booth_integrtaion_6_shift_reg_output_9, 
         booth_booth_integrtaion_6_shift_Reg_count_9, 
         booth_booth_integrtaion_6_shift_Reg_output_8, 
         booth_booth_integrtaion_6_shift_Reg_count_8, 
         booth_booth_integrtaion_6_shift_Reg_output_7, 
         booth_booth_integrtaion_6_shift_Reg_count_7, 
         booth_booth_integrtaion_6_shift_Reg_output_6, 
         booth_booth_integrtaion_6_shift_Reg_count_6, 
         booth_booth_integrtaion_6_shift_Reg_output_5, 
         booth_booth_integrtaion_6_shift_Reg_count_5, 
         booth_booth_integrtaion_6_shift_Reg_output_4, 
         booth_booth_integrtaion_6_shift_Reg_count_4, 
         booth_booth_integrtaion_6_shift_Reg_output_3, 
         booth_booth_integrtaion_6_shift_Reg_count_3, 
         booth_booth_integrtaion_6_shift_Reg_output_2, 
         booth_booth_integrtaion_6_shift_Reg_count_2, 
         booth_booth_integrtaion_6_shift_Reg_output_1, 
         booth_booth_integrtaion_6_shift_Reg_count_1, 
         booth_booth_integrtaion_6_shift_reg_output_0, 
         booth_booth_integrtaion_6_shift_Reg_count_0, 
         booth_booth_integration_output_6_1, booth_booth_integration_output_6_2, 
         booth_booth_integration_output_6_3, booth_booth_integration_output_6_4, 
         booth_booth_integration_output_6_5, booth_booth_integration_output_6_6, 
         booth_booth_integration_output_6_7, booth_booth_integration_output_6_8, 
         booth_booth_integration_output_6_9, booth_booth_integration_output_6_10, 
         booth_booth_integration_output_6_11, 
         booth_booth_integration_output_6_12, 
         booth_booth_integration_output_6_13, 
         booth_booth_integration_output_6_14, 
         booth_booth_integration_output_6_15, 
         booth_booth_integrtaion_6_booth_output_16, nx12836, nx12842, 
         booth_booth_integrtaion_6_booth_output_17, nx13296, nx12850, nx12866, 
         booth_booth_integrtaion_6_booth_output_18, nx13297, nx12876, nx12880, 
         nx12894, booth_booth_integrtaion_6_booth_output_19, nx13298, nx12900, 
         nx12904, nx12914, booth_booth_integrtaion_6_booth_output_20, nx13299, 
         nx12924, nx12928, nx12942, booth_booth_integrtaion_6_booth_output_21, 
         nx13300, nx12948, nx12952, nx12962, 
         booth_booth_integrtaion_6_booth_output_22, nx13301, nx12972, nx12976, 
         nx12990, booth_booth_integrtaion_6_booth_output_23, nx13303, nx12996, 
         nx13000, nx13010, booth_booth_integrtaion_6_booth_output_24, nx13305, 
         nx13020, nx13024, nx13038, booth_booth_integrtaion_6_booth_output_25, 
         nx13307, nx13044, nx13048, nx13058, 
         booth_booth_integrtaion_6_booth_output_26, nx13308, nx13068, nx13072, 
         nx13086, booth_booth_integrtaion_6_booth_output_27, nx13309, nx13092, 
         nx13096, nx13106, booth_booth_integrtaion_6_booth_output_28, nx13310, 
         nx13116, nx13120, nx13134, booth_booth_integrtaion_6_booth_output_29, 
         nx13311, nx13140, nx13144, nx13154, 
         booth_booth_integrtaion_6_booth_output_31, nx13312, nx13164, nx13168, 
         nx13182, nx13184, nx13192, nx13198, nx13206, nx13222, nx13230, nx13246, 
         nx13254, nx13270, nx13278, nx13294, nx13302, nx13318, nx13326, nx13342, 
         nx13350, nx13366, nx13372, nx13378, nx13396, nx13408, nx13420, nx13432, 
         nx13444, nx13456, nx13468, nx13480, nx13492, nx13504, nx13516, nx13528, 
         nx13540, nx13552, nx13564, nx13574, label_7_input_state_machine_0, 
         nx13586, label_7_input_1, label_7_input_state_machine_1, nx13315, 
         nx13608, nx13612, label_7_input_2, label_7_input_state_machine_2, 
         nx13640, nx13644, nx13662, label_7_input_3, 
         label_7_input_state_machine_3, nx13319, nx13672, nx13676, 
         label_7_input_4, label_7_input_state_machine_4, nx13704, nx13708, 
         nx13726, label_7_input_5, label_7_input_state_machine_5, nx13321, 
         nx13736, nx13740, label_7_input_6, label_7_input_state_machine_6, 
         nx13768, nx13772, nx13790, label_7_input_7, 
         label_7_input_state_machine_7, nx13323, nx13800, nx13804, 
         label_7_input_8, label_7_input_state_machine_8, nx13832, nx13836, 
         nx13854, label_7_input_9, label_7_input_state_machine_9, nx13325, 
         nx13864, nx13868, label_7_input_10, label_7_input_state_machine_10, 
         nx13896, nx13900, nx13918, label_7_input_11, 
         label_7_input_state_machine_11, nx13329, nx13928, nx13932, 
         label_7_input_12, label_7_input_state_machine_12, nx13960, nx13964, 
         nx13982, label_7_input_13, label_7_input_state_machine_13, nx13332, 
         nx13992, nx13996, nx14018, nx14022, label_8_input_14, 
         label_8_input_state_machine_14, label_8_input_0, 
         booth_booth_integrtaion_7_shift_reg_output_9, 
         booth_booth_integrtaion_7_shift_Reg_count_9, 
         booth_booth_integrtaion_7_shift_Reg_output_8, 
         booth_booth_integrtaion_7_shift_Reg_count_8, 
         booth_booth_integrtaion_7_shift_Reg_output_7, 
         booth_booth_integrtaion_7_shift_Reg_count_7, 
         booth_booth_integrtaion_7_shift_Reg_output_6, 
         booth_booth_integrtaion_7_shift_Reg_count_6, 
         booth_booth_integrtaion_7_shift_Reg_output_5, 
         booth_booth_integrtaion_7_shift_Reg_count_5, 
         booth_booth_integrtaion_7_shift_Reg_output_4, 
         booth_booth_integrtaion_7_shift_Reg_count_4, 
         booth_booth_integrtaion_7_shift_Reg_output_3, 
         booth_booth_integrtaion_7_shift_Reg_count_3, 
         booth_booth_integrtaion_7_shift_Reg_output_2, 
         booth_booth_integrtaion_7_shift_Reg_count_2, 
         booth_booth_integrtaion_7_shift_Reg_output_1, 
         booth_booth_integrtaion_7_shift_Reg_count_1, 
         booth_booth_integrtaion_7_shift_reg_output_0, 
         booth_booth_integrtaion_7_shift_Reg_count_0, 
         booth_booth_integration_output_7_1, booth_booth_integration_output_7_2, 
         booth_booth_integration_output_7_3, booth_booth_integration_output_7_4, 
         booth_booth_integration_output_7_5, booth_booth_integration_output_7_6, 
         booth_booth_integration_output_7_7, booth_booth_integration_output_7_8, 
         booth_booth_integration_output_7_9, booth_booth_integration_output_7_10, 
         booth_booth_integration_output_7_11, 
         booth_booth_integration_output_7_12, 
         booth_booth_integration_output_7_13, 
         booth_booth_integration_output_7_14, 
         booth_booth_integration_output_7_15, 
         booth_booth_integrtaion_7_booth_output_16, nx14152, nx14158, 
         booth_booth_integrtaion_7_booth_output_17, nx13334, nx14166, nx14182, 
         booth_booth_integrtaion_7_booth_output_18, nx13335, nx14192, nx14196, 
         nx14210, booth_booth_integrtaion_7_booth_output_19, nx13336, nx14216, 
         nx14220, nx14230, booth_booth_integrtaion_7_booth_output_20, nx13337, 
         nx14240, nx14244, nx14258, booth_booth_integrtaion_7_booth_output_21, 
         nx13339, nx14264, nx14268, nx14278, 
         booth_booth_integrtaion_7_booth_output_22, nx13341, nx14288, nx14292, 
         nx14306, booth_booth_integrtaion_7_booth_output_23, nx13343, nx14312, 
         nx14316, nx14326, booth_booth_integrtaion_7_booth_output_24, nx13344, 
         nx14336, nx14340, nx14354, booth_booth_integrtaion_7_booth_output_25, 
         nx13345, nx14360, nx14364, nx14374, 
         booth_booth_integrtaion_7_booth_output_26, nx13346, nx14384, nx14388, 
         nx14402, booth_booth_integrtaion_7_booth_output_27, nx13347, nx14408, 
         nx14412, nx14422, booth_booth_integrtaion_7_booth_output_28, nx13348, 
         nx14432, nx14436, nx14450, booth_booth_integrtaion_7_booth_output_29, 
         nx13349, nx14456, nx14460, nx14470, 
         booth_booth_integrtaion_7_booth_output_31, nx13351, nx14480, nx14484, 
         nx14498, nx14500, nx14508, nx14514, nx14522, nx14538, nx14546, nx14562, 
         nx14570, nx14586, nx14594, nx14610, nx14618, nx14634, nx14642, nx14658, 
         nx14666, nx14682, nx14688, nx14694, nx14712, nx14724, nx14736, nx14748, 
         nx14760, nx14772, nx14784, nx14796, nx14808, nx14820, nx14832, nx14844, 
         nx14856, nx14868, nx14880, nx14890, label_8_input_state_machine_0, 
         nx14902, label_8_input_1, label_8_input_state_machine_1, nx13355, 
         nx14924, nx14928, label_8_input_2, label_8_input_state_machine_2, 
         nx14956, nx14960, nx14978, label_8_input_3, 
         label_8_input_state_machine_3, nx13357, nx14988, nx14992, 
         label_8_input_4, label_8_input_state_machine_4, nx15020, nx15024, 
         nx15042, label_8_input_5, label_8_input_state_machine_5, nx13359, 
         nx15052, nx15056, label_8_input_6, label_8_input_state_machine_6, 
         nx15084, nx15088, nx15106, label_8_input_7, 
         label_8_input_state_machine_7, nx13361, nx15116, nx15120, 
         label_8_input_8, label_8_input_state_machine_8, nx15148, nx15152, 
         nx15170, label_8_input_9, label_8_input_state_machine_9, nx13365, 
         nx15180, nx15184, label_8_input_10, label_8_input_state_machine_10, 
         nx15212, nx15216, nx15234, label_8_input_11, 
         label_8_input_state_machine_11, nx13368, nx15244, nx15248, 
         label_8_input_12, label_8_input_state_machine_12, nx15276, nx15280, 
         nx15298, label_8_input_13, label_8_input_state_machine_13, nx13370, 
         nx15308, nx15312, nx15334, nx15338, nx15360, 
         max_calc_comparator_fourth_inp2_13, max_calc_comparator_fourth_inp1_13, 
         max_calc_comparator_fourth_inp1_12, nx15404, 
         max_calc_comparator_fourth_inp2_11, max_calc_comparator_fourth_inp1_11, 
         max_calc_comparator_fourth_inp1_10, nx15448, 
         max_calc_comparator_fourth_inp2_9, max_calc_comparator_fourth_inp1_9, 
         max_calc_comparator_fourth_inp1_8, nx15492, 
         max_calc_comparator_fourth_inp2_7, max_calc_comparator_fourth_inp1_7, 
         max_calc_comparator_fourth_inp1_6, nx15536, 
         max_calc_comparator_fourth_inp2_5, max_calc_comparator_fourth_inp1_5, 
         max_calc_comparator_fourth_inp1_4, nx15580, 
         max_calc_comparator_fourth_inp2_3, max_calc_comparator_fourth_inp1_3, 
         max_calc_comparator_fourth_inp1_2, nx15624, 
         max_calc_comparator_fourth_inp2_1, nx15646, 
         max_calc_comparator_fourth_inp1_0, nx15682, nx15698, nx15714, nx15730, 
         nx15746, nx15762, nx15778, label_8_input_15, 
         label_8_input_state_machine_15, nx15800, nx15804, nx15808, 
         label_7_input_15, label_7_input_state_machine_15, nx15842, nx15846, 
         nx15850, nx15872, nx15874, nx15896, nx15908, 
         max_calc_comparator_second_inp2_13, max_calc_ans4_13, nx15934, 
         max_calc_comparator_second_inp1_13, max_calc_ans3_13, nx15970, 
         max_calc_ans4_12, nx16008, max_calc_comparator_second_inp1_12, 
         max_calc_ans3_12, nx16044, nx16056, max_calc_comparator_second_inp2_11, 
         max_calc_ans4_11, nx16082, max_calc_comparator_second_inp1_11, 
         max_calc_ans3_11, nx16118, max_calc_ans4_10, nx16156, 
         max_calc_comparator_second_inp1_10, max_calc_ans3_10, nx16192, nx16204, 
         max_calc_comparator_second_inp2_9, max_calc_ans4_9, nx16230, 
         max_calc_comparator_second_inp1_9, max_calc_ans3_9, nx16266, 
         max_calc_ans4_8, nx16304, max_calc_comparator_second_inp1_8, 
         max_calc_ans3_8, nx16340, nx16352, max_calc_comparator_second_inp2_7, 
         max_calc_ans4_7, nx16378, max_calc_comparator_second_inp1_7, 
         max_calc_ans3_7, nx16414, max_calc_ans4_6, nx16452, 
         max_calc_comparator_second_inp1_6, max_calc_ans3_6, nx16488, nx16500, 
         max_calc_comparator_second_inp2_5, max_calc_ans4_5, nx16526, 
         max_calc_comparator_second_inp1_5, max_calc_ans3_5, nx16562, 
         max_calc_ans4_4, nx16600, max_calc_comparator_second_inp1_4, 
         max_calc_ans3_4, nx16636, nx16648, max_calc_comparator_second_inp2_3, 
         max_calc_ans4_3, nx16674, max_calc_comparator_second_inp1_3, 
         max_calc_ans3_3, nx16710, max_calc_ans4_2, nx16748, 
         max_calc_comparator_second_inp1_2, max_calc_ans3_2, nx16784, nx16796, 
         max_calc_comparator_second_inp2_1, max_calc_ans4_1, nx16822, 
         max_calc_ans3_1, nx16858, nx16870, max_calc_ans4_0, nx16896, 
         max_calc_comparator_second_inp1_0, max_calc_ans3_0, nx16932, nx16958, 
         nx16974, nx16990, nx17006, nx17022, nx17038, nx17054, max_calc_ans4_15, 
         nx17088, max_calc_ans3_15, nx17124, nx17136, nx17138, nx17146, nx17156, 
         max_calc_ans8_14, max_calc_comparator_first_inp1_14, max_calc_ans1_14, 
         nx13371, nx17174, max_calc_ans6_14, max_calc_ans5_14, nx17196, nx17206, 
         nx17210, nx13373, max_calc_ans7_14, nx17244, nx17248, nx17256, 
         max_calc_comparator_first_inp2_13, max_calc_ans2_13, nx17268, nx17278, 
         max_calc_ans8_13, max_calc_comparator_first_inp1_13, max_calc_ans1_13, 
         nx13375, nx17296, max_calc_ans6_13, max_calc_ans5_13, nx17318, nx17328, 
         nx17332, max_calc_ans7_13, nx17366, nx17370, 
         max_calc_comparator_first_inp2_12, max_calc_ans2_12, nx17390, nx17400, 
         max_calc_ans8_12, max_calc_comparator_first_inp1_12, max_calc_ans1_12, 
         nx13376, nx17418, max_calc_ans6_12, max_calc_ans5_12, nx17440, nx17450, 
         nx17454, max_calc_ans7_12, nx17488, nx17492, nx17500, 
         max_calc_comparator_first_inp2_11, max_calc_ans2_11, nx17512, nx17522, 
         max_calc_ans8_11, max_calc_comparator_first_inp1_11, max_calc_ans1_11, 
         nx13377, nx17540, max_calc_ans6_11, max_calc_ans5_11, nx17562, nx17572, 
         nx17576, max_calc_ans7_11, nx17610, nx17614, 
         max_calc_comparator_first_inp2_10, max_calc_ans2_10, nx17634, nx17644, 
         max_calc_ans8_10, max_calc_comparator_first_inp1_10, max_calc_ans1_10, 
         nx13379, nx17662, max_calc_ans6_10, max_calc_ans5_10, nx17684, nx17694, 
         nx17698, max_calc_ans7_10, nx17732, nx17736, nx17744, 
         max_calc_comparator_first_inp2_9, max_calc_ans2_9, nx17756, nx17766, 
         max_calc_ans8_9, max_calc_comparator_first_inp1_9, max_calc_ans1_9, 
         nx13381, nx17784, max_calc_ans6_9, max_calc_ans5_9, nx17806, nx17816, 
         nx17820, max_calc_ans7_9, nx17854, nx17858, 
         max_calc_comparator_first_inp2_8, max_calc_ans2_8, nx17878, nx17888, 
         max_calc_ans8_8, max_calc_comparator_first_inp1_8, max_calc_ans1_8, 
         nx13383, nx17906, max_calc_ans6_8, max_calc_ans5_8, nx17928, nx17938, 
         nx17942, max_calc_ans7_8, nx17976, nx17980, nx17988, 
         max_calc_comparator_first_inp2_7, max_calc_ans2_7, nx18000, nx18010, 
         max_calc_ans8_7, max_calc_comparator_first_inp1_7, max_calc_ans1_7, 
         nx13385, nx18028, max_calc_ans6_7, max_calc_ans5_7, nx18050, nx18060, 
         nx18064, max_calc_ans7_7, nx18098, nx18102, 
         max_calc_comparator_first_inp2_6, max_calc_ans2_6, nx18122, nx18132, 
         max_calc_ans8_6, max_calc_comparator_first_inp1_6, max_calc_ans1_6, 
         nx13386, nx18150, max_calc_ans6_6, max_calc_ans5_6, nx18172, nx18182, 
         nx18186, max_calc_ans7_6, nx18220, nx18224, nx18232, 
         max_calc_comparator_first_inp2_5, max_calc_ans2_5, nx18244, nx18254, 
         max_calc_ans8_5, max_calc_comparator_first_inp1_5, max_calc_ans1_5, 
         nx13387, nx18272, max_calc_ans6_5, max_calc_ans5_5, nx18294, nx18304, 
         nx18308, max_calc_ans7_5, nx18342, nx18346, 
         max_calc_comparator_first_inp2_4, max_calc_ans2_4, nx18366, nx18376, 
         max_calc_ans8_4, max_calc_comparator_first_inp1_4, max_calc_ans1_4, 
         nx13388, nx18394, max_calc_ans6_4, max_calc_ans5_4, nx18416, nx18426, 
         nx18430, max_calc_ans7_4, nx18464, nx18468, nx18476, 
         max_calc_comparator_first_inp2_3, max_calc_ans2_3, nx18488, nx18498, 
         max_calc_ans8_3, max_calc_comparator_first_inp1_3, max_calc_ans1_3, 
         nx13389, nx18516, max_calc_ans6_3, max_calc_ans5_3, nx18538, nx18548, 
         nx18552, max_calc_ans7_3, nx18586, nx18590, 
         max_calc_comparator_first_inp2_2, max_calc_ans2_2, nx18610, nx18620, 
         max_calc_ans8_2, max_calc_comparator_first_inp1_2, max_calc_ans1_2, 
         nx13391, nx18638, max_calc_ans6_2, max_calc_ans5_2, nx18660, nx18670, 
         nx18674, max_calc_ans7_2, nx18708, nx18712, nx18720, 
         max_calc_comparator_first_inp2_1, max_calc_ans2_1, nx18732, nx18742, 
         max_calc_ans8_1, max_calc_comparator_first_inp1_1, max_calc_ans1_1, 
         nx13393, nx18760, max_calc_ans6_1, max_calc_ans5_1, nx18782, nx18792, 
         nx18796, max_calc_ans7_1, nx18830, nx18834, nx18842, 
         max_calc_comparator_first_inp2_0, max_calc_ans2_0, nx18854, nx18864, 
         max_calc_ans8_0, max_calc_ans7_0, nx18888, nx18892, nx18914, nx18930, 
         nx18946, nx18962, nx18978, nx18994, nx19010, 
         max_calc_comparator_first_inp2_15, max_calc_ans2_15, nx19030, nx19040, 
         max_calc_ans8_15, max_calc_comparator_first_inp1_15, max_calc_ans1_15, 
         nx13395, nx19058, max_calc_ans6_15, max_calc_ans5_15, nx19080, nx19090, 
         nx19094, max_calc_ans7_15, nx19128, nx19132, nx19140, nx19232, nx19236, 
         nx19240, nx19250, nx19266, nx19276, nx19296, nx13403, nx13413, nx13423, 
         nx13429, nx13443, nx13453, nx13463, nx13473, nx13483, nx13493, nx13503, 
         nx13513, nx13523, nx13533, nx13543, nx13553, nx13563, nx13573, nx13583, 
         nx13593, nx13603, nx13613, nx13623, nx13633, nx13643, nx13653, nx13663, 
         nx13673, nx13683, nx13693, nx13703, nx13713, nx13723, nx13733, nx13743, 
         nx13753, nx13763, nx13773, nx13783, nx13793, nx13803, nx13813, nx13823, 
         nx13833, nx13843, nx13853, nx13863, nx13873, nx13883, nx13893, nx13903, 
         nx13913, nx13923, nx13933, nx13943, nx13953, nx13963, nx13973, nx13983, 
         nx13993, nx14003, nx14013, nx14023, nx14033, nx14043, nx14053, nx14063, 
         nx14073, nx14083, nx14093, nx14103, nx14113, nx14123, nx14133, nx14139, 
         nx14153, nx14163, nx14173, nx14183, nx14193, nx14203, nx14213, nx14223, 
         nx14233, nx14243, nx14253, nx14263, nx14273, nx14283, nx14293, nx14303, 
         nx14313, nx14323, nx14333, nx14343, nx14353, nx14363, nx14373, nx14383, 
         nx14393, nx14403, nx14413, nx14423, nx14433, nx14443, nx14453, nx14463, 
         nx14473, nx14483, nx14493, nx14503, nx14513, nx14523, nx14533, nx14543, 
         nx14553, nx14563, nx14573, nx14583, nx14593, nx14603, nx14613, nx14623, 
         nx14633, nx14643, nx14653, nx14663, nx14673, nx14683, nx14693, nx14703, 
         nx14713, nx14723, nx14733, nx14743, nx14753, nx14763, nx14773, nx14783, 
         nx14793, nx14803, nx14813, nx14823, nx14833, nx14843, nx14853, nx14863, 
         nx14873, nx14883, nx14893, nx14903, nx14913, nx14923, nx14933, nx14943, 
         nx14953, nx14963, nx14973, nx14983, nx14989, nx15003, nx15013, nx15023, 
         nx15033, nx15043, nx15053, nx15063, nx15073, nx15083, nx15093, nx15103, 
         nx15113, nx15123, nx15133, nx15143, nx15153, nx15163, nx15173, nx15183, 
         nx15193, nx15203, nx15213, nx15223, nx15233, nx15243, nx15253, nx15263, 
         nx15273, nx15283, nx15293, nx15303, nx15313, nx15323, nx15333, nx15343, 
         nx15353, nx15363, nx15373, nx15383, nx15393, nx15403, nx15413, nx15423, 
         nx15433, nx15443, nx15453, nx15463, nx15473, nx15483, nx15493, nx15503, 
         nx15513, nx15523, nx15533, nx15543, nx15553, nx15563, nx15573, nx15583, 
         nx15593, nx15603, nx15613, nx15623, nx15633, nx15643, nx15653, nx15663, 
         nx15673, nx15683, nx15693, nx15703, nx15713, nx15723, nx15733, nx15743, 
         nx15753, nx15763, nx15773, nx15783, nx15793, nx15803, nx15813, nx15823, 
         nx15833, nx15839, nx15853, nx15863, nx15873, nx15883, nx15893, nx15903, 
         nx15913, nx15923, nx15933, nx15943, nx15953, nx15963, nx15973, nx15983, 
         nx15993, nx16003, nx16013, nx16023, nx16033, nx16043, nx16053, nx16063, 
         nx16073, nx16083, nx16093, nx16103, nx16113, nx16123, nx16133, nx16143, 
         nx16153, nx16163, nx16173, nx16183, nx16193, nx16203, nx16213, nx16223, 
         nx16233, nx16243, nx16253, nx16263, nx16273, nx16283, nx16293, nx16303, 
         nx16313, nx16323, nx16333, nx16343, nx16353, nx16363, nx16373, nx16383, 
         nx16393, nx16403, nx16413, nx16423, nx16433, nx16443, nx16453, nx16463, 
         nx16473, nx16483, nx16493, nx16503, nx16513, nx16523, nx16533, nx16543, 
         nx16553, nx16563, nx16573, nx16583, nx16593, nx16603, nx16613, nx16623, 
         nx16633, nx16643, nx16653, nx16663, nx16673, nx16683, nx16689, nx16703, 
         nx16713, nx16723, nx16733, nx16743, nx16753, nx16763, nx16773, nx16783, 
         nx16793, nx16803, nx16813, nx16823, nx16833, nx16843, nx16853, nx16863, 
         nx16873, nx16883, nx16893, nx16903, nx16913, nx16923, nx16933, nx16943, 
         nx16953, nx16963, nx16973, nx16983, nx16993, nx17003, nx17013, nx17023, 
         nx17033, nx17043, nx17053, nx17063, nx17073, nx17083, nx17093, nx17103, 
         nx17113, nx17123, nx17133, nx17143, nx17153, nx17163, nx17173, nx17183, 
         nx17193, nx17203, nx17213, nx17223, nx17233, nx17243, nx17253, nx17263, 
         nx17273, nx17283, nx17293, nx17303, nx17313, nx17323, nx17333, nx17343, 
         nx17353, nx17363, nx17373, nx17383, nx17393, nx17403, nx17413, nx17423, 
         nx17433, nx17443, nx17453, nx17463, nx17473, nx17483, nx17493, nx17503, 
         nx17513, nx17523, nx17533, nx17543, nx17553, nx17563, nx17573, nx17583, 
         nx17593, nx17603, nx17609, nx17623, nx17633, nx17643, nx17653, nx17663, 
         nx17673, nx17683, nx17693, nx17703, nx17713, nx17723, nx17733, nx17743, 
         nx17753, nx17763, nx17773, nx17783, nx17793, nx17803, nx17813, nx17823, 
         nx17833, nx17843, nx17853, nx17863, nx17873, nx17883, nx17893, nx17903, 
         nx17913, nx17923, nx17933, nx17943, nx17953, nx17963, nx17973, nx17983, 
         nx17993, nx18003, nx18013, nx18023, nx18033, nx18043, nx18053, nx18063, 
         nx18073, nx18083, nx18093, nx18103, nx18113, nx18123, nx18133, nx18143, 
         nx18153, nx18163, nx18173, nx18179, nx18193, nx18203, nx18213, nx18223, 
         nx18233, nx18243, nx18253, nx18263, nx18273, nx18283, nx18293, nx18303, 
         nx18313, nx18323, nx18333, nx18343, nx18353, nx18363, nx18373, nx18383, 
         nx18393, nx18403, nx18413, nx18423, nx18433, nx18443, nx18453, nx18463, 
         nx18473, nx18483, nx18493, nx18503, nx18513, nx18523, nx18533, nx18543, 
         nx18553, nx18563, nx18573, nx18583, nx18593, nx18603, nx18613, nx18623, 
         nx18633, nx18643, nx18653, nx18663, nx18673, nx18683, nx18693, nx18703, 
         nx18713, nx18723, nx18733, nx18743, nx18753, nx18763, nx18773, nx18783, 
         nx18793, nx18803, nx18813, nx18823, nx18833, nx18843, nx18853, nx18863, 
         nx18873, nx18883, nx18893, nx18903, nx18913, nx18923, nx18933, nx18943, 
         nx18953, nx18963, nx18973, nx18983, nx18993, nx19003, nx19013, nx19023, 
         nx19033, nx19043, nx19053, nx19063, nx19073, nx19083, nx19093, nx19103, 
         nx19113, nx19123, nx19133, nx19143, nx19153, nx19163, nx19173, nx19183, 
         nx19193, nx19203, nx19213, nx19223, nx19233, nx19243, nx19253, nx19263, 
         nx19273, nx19283, nx19293, nx19303, nx19313, nx19323, nx19333, nx19343, 
         nx19353, nx19363, nx19373, nx19383, nx19393, nx19403, nx19413, nx19423, 
         nx19433, nx19443, nx19453, nx19463, nx19473, nx19483, nx19493, nx19503, 
         nx19513, nx19523, nx19533, nx19543, nx19553, nx19563, nx19573, nx19583, 
         nx19593, nx19603, nx19613, nx19623, nx19633, nx19643, nx19653, nx19659, 
         nx19673, nx19683, nx19693, nx19703, nx19713, nx19723, nx19733, nx19743, 
         nx19753, nx19763, nx19773, nx19783, nx19793, nx19803, nx19813, nx19823, 
         nx19833, nx19843, nx19853, nx19863, nx19873, nx19883, nx19893, nx19903, 
         nx19913, nx19923, nx19933, nx19943, nx19953, nx19963, nx19973, nx19983, 
         nx19993, nx20003, nx20013, nx20023, nx20033, nx20043, nx20053, nx20063, 
         nx20073, nx20083, nx20093, nx20103, nx20113, nx20123, nx20133, nx20143, 
         nx20153, nx20163, nx20173, nx20183, nx20193, nx20203, nx20213, nx20223, 
         nx20233, nx20243, nx20253, nx20263, nx20273, nx20283, nx20293, nx20303, 
         nx20313, nx20323, nx20333, nx20343, nx20353, nx20363, nx20373, nx20383, 
         nx20393, nx20403, nx20413, nx20423, nx20433, nx20443, nx20453, nx20463, 
         nx20473, nx20483, nx20493, nx20499, nx20513, nx20523, nx20533, nx20543, 
         nx20553, nx20563, nx20573, nx20583, nx20593, nx20603, nx20613, nx20623, 
         nx20633, nx20643, nx20653, nx20663, nx20673, nx20683, nx20693, nx20703, 
         nx20713, nx20723, nx20733, nx20743, nx20753, nx20763, nx20773, nx20783, 
         nx20793, nx20803, nx20813, nx20823, nx20833, nx20843, nx20853, nx20863, 
         nx20873, nx20883, nx20893, nx20903, nx20913, nx20923, nx20933, nx20943, 
         nx20953, nx20963, nx20973, nx20983, nx20993, nx21003, nx21013, nx21023, 
         nx21033, nx21043, nx21053, nx21063, nx21073, nx21083, nx21093, nx21103, 
         nx21113, nx21123, nx21133, nx21143, nx21153, nx21163, nx21173, nx21183, 
         nx21193, nx21203, nx21213, nx21223, nx21233, nx21243, nx21253, nx21263, 
         nx21273, nx21283, nx21293, nx21303, nx21313, nx21323, nx21333, nx21343, 
         nx21353, nx21363, nx21373, nx21383, nx21393, nx21403, nx21413, nx21423, 
         nx21433, nx21443, nx21453, nx21463, nx21473, nx21483, nx21493, nx21503, 
         nx21513, nx21523, nx21533, nx21543, nx21553, nx21563, nx21573, nx21583, 
         nx21593, nx21603, nx21613, nx21623, nx21633, nx21643, nx21653, nx21663, 
         nx21673, nx21683, nx21693, nx21699, nx21713, nx21723, nx21733, nx21743, 
         nx21753, nx21763, nx21773, nx21783, nx21793, nx21803, nx21813, nx21823, 
         nx21833, nx21843, nx21853, nx21863, nx21873, nx21883, nx21893, nx21903, 
         nx21913, nx21923, nx21933, nx21943, nx21953, nx21963, nx21973, nx21983, 
         nx21993, nx22003, nx22013, nx22023, nx22033, nx22043, nx22053, nx22063, 
         nx22073, nx22083, nx22093, nx22103, nx22113, nx22123, nx22133, nx22143, 
         nx22153, nx22163, nx22173, nx22183, nx22193, nx22203, nx22213, nx22223, 
         nx22233, nx22243, nx22253, nx22263, nx22273, nx22283, nx22293, nx22303, 
         nx22313, nx22323, nx22333, nx22343, nx22353, nx22363, nx22373, nx22383, 
         nx22393, nx22403, nx22413, nx22423, nx22433, nx22443, nx22453, nx22463, 
         nx22473, nx22483, nx22493, nx22503, nx22513, nx22523, nx22533, nx22539, 
         nx22553, nx22563, nx22573, nx22583, nx22593, nx22603, nx22613, nx22623, 
         nx22633, nx22643, nx22653, nx22663, nx22673, nx22683, nx22693, nx22703, 
         nx22713, nx22723, nx22733, nx22743, nx22753, nx22763, nx22773, nx22783, 
         nx22793, nx22803, nx22813, nx22823, nx22833, nx22843, nx22853, nx22863, 
         nx22873, nx22883, nx22893, nx22903, nx22913, nx22923, nx22933, nx22943, 
         nx22953, nx22963, nx22973, nx22983, nx22993, nx23003, nx23013, nx23023, 
         nx23033, nx23043, nx23053, nx23063, nx23073, nx23083, nx23093, nx23103, 
         nx23113, nx23123, nx23133, nx23143, nx23153, nx23163, nx23173, nx23183, 
         nx23193, nx23203, nx23213, nx23223, nx23233, nx23243, nx23253, nx23263, 
         nx23273, nx23283, nx23293, nx23303, nx23313, nx23323, nx23333, nx23343, 
         nx23353, nx23363, nx23373, nx23383, nx23393, nx23403, nx23413, nx23423, 
         nx23433, nx23443, nx23453, nx23463, nx23473, nx23483, nx23493, nx23503, 
         nx23513, nx23523, nx23533, nx23543, nx23553, nx23563, nx23573, nx23583, 
         nx23593, nx23603, nx23613, nx23623, nx23633, nx23643, nx23653, nx23663, 
         nx23673, nx23683, nx23693, nx23703, nx23713, nx23723, nx23733, nx23743, 
         nx23753, nx23763, nx23773, nx23783, nx23793, nx23803, nx23813, nx23823, 
         nx23833, nx23843, nx23853, nx23863, nx23873, nx23883, nx23893, nx23903, 
         nx23913, nx23923, nx23933, nx23943, nx23953, nx23963, nx23973, nx23983, 
         nx23993, nx24003, nx24013, nx24023, nx24033, nx24043, nx24053, nx24063, 
         nx24073, nx24083, nx24093, nx24103, nx24113, nx24123, nx24133, nx24143, 
         nx24153, nx24163, nx24173, nx24183, nx24193, nx24203, nx24213, nx24223, 
         nx24233, nx24243, nx24253, nx24263, nx24273, nx24283, nx24293, nx24303, 
         nx24313, nx24323, nx24333, nx24343, nx24353, nx24363, nx24373, nx24383, 
         nx24393, nx24403, nx24413, nx24423, nx24433, nx24443, nx24453, nx24463, 
         nx24473, nx24483, nx24493, nx24503, nx24513, nx24523, nx24533, nx24543, 
         nx24553, nx24563, nx24573, nx24583, nx24593, nx24603, nx24613, nx24623, 
         nx24633, nx24643, nx24653, nx24663, nx24673, nx24683, nx24693, nx24703, 
         nx24713, nx24723, nx24733, nx24743, nx24753, nx24763, nx24773, nx24783, 
         nx24793, nx24803, nx24813, nx24823, nx24833, nx24843, nx24853, nx24863, 
         nx24873, nx24883, nx24893, nx24903, nx24913, nx24923, nx24933, nx24943, 
         nx24953, nx24963, nx24973, nx24983, nx24993, nx25003, nx25013, nx25023, 
         nx25033, nx25043, nx25053, nx25063, nx25073, nx25083, nx25093, nx25103, 
         nx25113, nx25123, nx25133, nx25143, nx25153, nx25163, nx25173, nx25183, 
         nx25193, nx25203, nx25213, nx25223, nx25233, nx25243, nx25253, nx25263, 
         nx25273, nx25283, nx25293, nx25303, nx25313, nx25323, nx25333, nx25343, 
         nx25353, nx25363, nx25373, nx25383, nx25393, nx25403, nx25413, nx25423, 
         nx25433, nx25443, nx25453, nx25463, nx25473, nx25483, nx25493, nx25503, 
         nx25513, nx25523, nx25533, nx25543, nx25553, nx25563, nx25573, nx25583, 
         nx25593, nx25603, nx25613, nx25623, nx25633, nx25643, nx25653, nx25663, 
         nx25673, nx25683, nx25693, nx25703, nx25713, nx25723, nx25733, nx25743, 
         nx25753, nx25757, nx25813, nx25821, nx25823, nx25827, nx25830, nx25832, 
         nx25835, nx25849, nx25854, nx25857, nx25864, nx25874, nx25879, nx25891, 
         nx25893, nx25896, nx25900, nx25902, nx25907, nx25916, nx25919, nx25935, 
         nx25937, nx25940, nx25942, nx25944, nx25949, nx25951, nx25958, nx25962, 
         nx25975, nx25982, nx25986, nx25998, nx25999, nx26001, nx26014, nx26022, 
         nx26024, nx26027, nx26039, nx26044, nx26046, nx26052, nx26056, nx26069, 
         nx26078, nx26080, nx26083, nx26095, nx26099, nx26105, nx26109, nx26122, 
         nx26129, nx26144, nx26176, nx26180, nx26182, nx26184, nx26186, nx26188, 
         nx26191, nx26194, nx26201, nx26203, nx26223, nx26227, nx26276, nx26323, 
         nx26344, nx26349, nx26351, nx26353, nx26356, nx26360, nx26366, nx26368, 
         nx26371, nx26375, nx26381, nx26384, nx26386, nx26389, nx26391, nx26396, 
         nx26398, nx26401, nx26404, nx26412, nx26418, nx26421, nx26423, nx26426, 
         nx26428, nx26430, nx26435, nx26437, nx26440, nx26443, nx26453, nx26456, 
         nx26458, nx26461, nx26463, nx26465, nx26470, nx26472, nx26475, nx26478, 
         nx26488, nx26491, nx26493, nx26496, nx26498, nx26500, nx26505, nx26507, 
         nx26510, nx26513, nx26523, nx26526, nx26528, nx26531, nx26533, nx26535, 
         nx26540, nx26542, nx26545, nx26548, nx26558, nx26561, nx26563, nx26566, 
         nx26568, nx26570, nx26575, nx26577, nx26580, nx26583, nx26593, nx26596, 
         nx26598, nx26601, nx26603, nx26605, nx26608, nx26612, nx26615, nx26618, 
         nx26621, nx26624, nx26627, nx26630, nx26634, nx26636, nx26638, nx26640, 
         nx26642, nx26644, nx26646, nx26648, nx26661, nx26664, nx26666, nx26669, 
         nx26675, nx26693, nx26696, nx26702, nx26706, nx26755, nx26802, nx26823, 
         nx26828, nx26830, nx26832, nx26835, nx26839, nx26845, nx26847, nx26850, 
         nx26854, nx26860, nx26863, nx26865, nx26868, nx26870, nx26875, nx26877, 
         nx26880, nx26883, nx26891, nx26897, nx26900, nx26902, nx26905, nx26907, 
         nx26909, nx26914, nx26916, nx26919, nx26922, nx26932, nx26935, nx26937, 
         nx26940, nx26942, nx26944, nx26949, nx26951, nx26954, nx26957, nx26967, 
         nx26970, nx26972, nx26975, nx26977, nx26979, nx26984, nx26986, nx26989, 
         nx26992, nx27002, nx27005, nx27007, nx27010, nx27012, nx27014, nx27019, 
         nx27021, nx27024, nx27027, nx27037, nx27040, nx27042, nx27045, nx27047, 
         nx27049, nx27054, nx27056, nx27059, nx27062, nx27072, nx27075, nx27077, 
         nx27080, nx27082, nx27084, nx27087, nx27091, nx27094, nx27097, nx27100, 
         nx27103, nx27106, nx27109, nx27113, nx27115, nx27117, nx27119, nx27121, 
         nx27123, nx27125, nx27127, nx27133, nx27135, nx27141, nx27145, nx27194, 
         nx27241, nx27262, nx27267, nx27269, nx27271, nx27274, nx27278, nx27284, 
         nx27286, nx27289, nx27293, nx27299, nx27302, nx27304, nx27307, nx27309, 
         nx27314, nx27316, nx27319, nx27322, nx27330, nx27336, nx27339, nx27341, 
         nx27344, nx27346, nx27348, nx27353, nx27355, nx27358, nx27361, nx27371, 
         nx27374, nx27376, nx27379, nx27381, nx27383, nx27388, nx27390, nx27393, 
         nx27396, nx27406, nx27409, nx27411, nx27414, nx27416, nx27418, nx27423, 
         nx27425, nx27428, nx27431, nx27441, nx27444, nx27446, nx27449, nx27451, 
         nx27453, nx27458, nx27460, nx27463, nx27466, nx27476, nx27479, nx27481, 
         nx27484, nx27486, nx27488, nx27493, nx27495, nx27498, nx27501, nx27511, 
         nx27514, nx27516, nx27519, nx27521, nx27523, nx27526, nx27530, nx27533, 
         nx27536, nx27539, nx27542, nx27545, nx27548, nx27552, nx27554, nx27556, 
         nx27558, nx27560, nx27562, nx27564, nx27566, nx27571, nx27573, nx27576, 
         nx27586, nx27597, nx27608, nx27619, nx27630, nx27641, nx27652, nx27663, 
         nx27665, nx27668, nx27678, nx27679, nx27683, nx27693, nx27694, nx27698, 
         nx27708, nx27709, nx27713, nx27723, nx27724, nx27728, nx27738, nx27739, 
         nx27743, nx27753, nx27754, nx27758, nx27760, nx27763, nx27765, nx27775, 
         nx27786, nx27797, nx27808, nx27819, nx27830, nx27841, nx27852, nx27854, 
         nx27857, nx27867, nx27868, nx27872, nx27882, nx27883, nx27887, nx27897, 
         nx27898, nx27902, nx27912, nx27913, nx27917, nx27927, nx27928, nx27932, 
         nx27942, nx27943, nx27947, nx27949, nx27952, nx27956, nx27958, nx27960, 
         nx27963, nx27965, nx27967, nx27970, nx27974, nx27976, nx27980, nx27984, 
         nx27986, nx27988, nx27991, nx27993, nx27995, nx27998, nx28002, nx28004, 
         nx28008, nx28012, nx28014, nx28016, nx28019, nx28021, nx28023, nx28026, 
         nx28030, nx28032, nx28036, nx28040, nx28042, nx28044, nx28047, nx28049, 
         nx28051, nx28054, nx28058, nx28060, nx28064, nx28068, nx28070, nx28072, 
         nx28075, nx28077, nx28079, nx28082, nx28086, nx28088, nx28092, nx28096, 
         nx28098, nx28100, nx28103, nx28105, nx28107, nx28110, nx28114, nx28116, 
         nx28122, nx28124, nx28126, nx28129, nx28131, nx28137, nx28139, nx28150, 
         nx28155, nx28157, nx28168, nx28172, nx28183, nx28187, nx28236, nx28283, 
         nx28304, nx28309, nx28311, nx28313, nx28316, nx28320, nx28326, nx28328, 
         nx28331, nx28335, nx28341, nx28344, nx28346, nx28349, nx28351, nx28356, 
         nx28358, nx28361, nx28364, nx28372, nx28378, nx28381, nx28383, nx28386, 
         nx28388, nx28390, nx28395, nx28397, nx28400, nx28403, nx28413, nx28416, 
         nx28418, nx28421, nx28423, nx28425, nx28430, nx28432, nx28435, nx28438, 
         nx28448, nx28451, nx28453, nx28456, nx28458, nx28460, nx28465, nx28467, 
         nx28470, nx28473, nx28483, nx28486, nx28488, nx28491, nx28493, nx28495, 
         nx28500, nx28502, nx28505, nx28508, nx28518, nx28521, nx28523, nx28526, 
         nx28528, nx28530, nx28535, nx28537, nx28540, nx28543, nx28553, nx28556, 
         nx28558, nx28561, nx28563, nx28565, nx28568, nx28572, nx28575, nx28578, 
         nx28581, nx28584, nx28587, nx28590, nx28594, nx28596, nx28598, nx28600, 
         nx28602, nx28604, nx28606, nx28608, nx28617, nx28619, nx28626, nx28630, 
         nx28679, nx28726, nx28747, nx28752, nx28754, nx28756, nx28759, nx28763, 
         nx28769, nx28771, nx28774, nx28778, nx28784, nx28787, nx28789, nx28792, 
         nx28794, nx28799, nx28801, nx28804, nx28807, nx28815, nx28821, nx28824, 
         nx28826, nx28829, nx28831, nx28833, nx28838, nx28840, nx28843, nx28846, 
         nx28856, nx28859, nx28861, nx28864, nx28866, nx28868, nx28873, nx28875, 
         nx28878, nx28881, nx28891, nx28894, nx28896, nx28899, nx28901, nx28903, 
         nx28908, nx28910, nx28913, nx28916, nx28926, nx28929, nx28931, nx28934, 
         nx28936, nx28938, nx28943, nx28945, nx28948, nx28951, nx28961, nx28964, 
         nx28966, nx28969, nx28971, nx28973, nx28978, nx28980, nx28983, nx28986, 
         nx28996, nx28999, nx29001, nx29004, nx29006, nx29008, nx29011, nx29015, 
         nx29018, nx29021, nx29024, nx29027, nx29030, nx29033, nx29037, nx29039, 
         nx29041, nx29043, nx29045, nx29047, nx29049, nx29051, nx29061, nx29063, 
         nx29069, nx29073, nx29122, nx29169, nx29190, nx29195, nx29197, nx29199, 
         nx29202, nx29206, nx29212, nx29214, nx29217, nx29221, nx29227, nx29230, 
         nx29232, nx29235, nx29237, nx29242, nx29244, nx29247, nx29250, nx29258, 
         nx29264, nx29267, nx29269, nx29272, nx29274, nx29276, nx29281, nx29283, 
         nx29286, nx29289, nx29299, nx29302, nx29304, nx29307, nx29309, nx29311, 
         nx29316, nx29318, nx29321, nx29324, nx29334, nx29337, nx29339, nx29342, 
         nx29344, nx29346, nx29351, nx29353, nx29356, nx29359, nx29369, nx29372, 
         nx29374, nx29377, nx29379, nx29381, nx29386, nx29388, nx29391, nx29394, 
         nx29404, nx29407, nx29409, nx29412, nx29414, nx29416, nx29421, nx29423, 
         nx29426, nx29429, nx29439, nx29442, nx29444, nx29447, nx29449, nx29451, 
         nx29454, nx29458, nx29461, nx29464, nx29467, nx29470, nx29473, nx29476, 
         nx29480, nx29482, nx29484, nx29486, nx29488, nx29490, nx29492, nx29494, 
         nx29498, nx29502, nx29504, nx29510, nx29514, nx29563, nx29610, nx29631, 
         nx29636, nx29638, nx29640, nx29643, nx29647, nx29653, nx29655, nx29658, 
         nx29662, nx29668, nx29671, nx29673, nx29676, nx29678, nx29683, nx29685, 
         nx29688, nx29691, nx29699, nx29705, nx29708, nx29710, nx29713, nx29715, 
         nx29717, nx29722, nx29724, nx29727, nx29730, nx29740, nx29743, nx29745, 
         nx29748, nx29750, nx29752, nx29757, nx29759, nx29762, nx29765, nx29775, 
         nx29778, nx29780, nx29783, nx29785, nx29787, nx29792, nx29794, nx29797, 
         nx29800, nx29810, nx29813, nx29815, nx29818, nx29820, nx29822, nx29827, 
         nx29829, nx29832, nx29835, nx29845, nx29848, nx29850, nx29853, nx29855, 
         nx29857, nx29862, nx29864, nx29867, nx29870, nx29880, nx29883, nx29885, 
         nx29888, nx29890, nx29892, nx29895, nx29899, nx29902, nx29905, nx29908, 
         nx29911, nx29914, nx29917, nx29921, nx29923, nx29925, nx29927, nx29929, 
         nx29931, nx29933, nx29935, nx29940, nx29942, nx29945, nx29955, nx29966, 
         nx29977, nx29988, nx29999, nx30010, nx30021, nx30032, nx30034, nx30037, 
         nx30047, nx30048, nx30052, nx30062, nx30063, nx30067, nx30077, nx30078, 
         nx30082, nx30092, nx30093, nx30097, nx30107, nx30108, nx30112, nx30122, 
         nx30123, nx30127, nx30129, nx30132, nx30134, nx30144, nx30155, nx30166, 
         nx30177, nx30188, nx30199, nx30210, nx30221, nx30223, nx30226, nx30236, 
         nx30237, nx30241, nx30251, nx30252, nx30256, nx30266, nx30267, nx30271, 
         nx30281, nx30282, nx30286, nx30296, nx30297, nx30301, nx30311, nx30312, 
         nx30316, nx30318, nx30321, nx30325, nx30327, nx30329, nx30332, nx30334, 
         nx30336, nx30339, nx30343, nx30345, nx30349, nx30353, nx30355, nx30357, 
         nx30360, nx30362, nx30364, nx30367, nx30371, nx30373, nx30377, nx30381, 
         nx30383, nx30385, nx30388, nx30390, nx30392, nx30395, nx30399, nx30401, 
         nx30405, nx30409, nx30411, nx30413, nx30416, nx30418, nx30420, nx30423, 
         nx30427, nx30429, nx30433, nx30437, nx30439, nx30441, nx30444, nx30446, 
         nx30448, nx30451, nx30455, nx30457, nx30461, nx30465, nx30467, nx30469, 
         nx30472, nx30474, nx30476, nx30479, nx30483, nx30485, nx30491, nx30493, 
         nx30495, nx30498, nx30500, nx30506, nx30508, nx30519, nx30524, nx30526, 
         nx30537, nx30546, nx30548, nx30555, nx30559, nx30608, nx30655, nx30676, 
         nx30681, nx30683, nx30685, nx30688, nx30692, nx30698, nx30700, nx30703, 
         nx30707, nx30713, nx30716, nx30718, nx30721, nx30723, nx30728, nx30730, 
         nx30733, nx30736, nx30744, nx30750, nx30753, nx30755, nx30758, nx30760, 
         nx30762, nx30767, nx30769, nx30772, nx30775, nx30785, nx30788, nx30790, 
         nx30793, nx30795, nx30797, nx30802, nx30804, nx30807, nx30810, nx30820, 
         nx30823, nx30825, nx30828, nx30830, nx30832, nx30837, nx30839, nx30842, 
         nx30845, nx30855, nx30858, nx30860, nx30863, nx30865, nx30867, nx30872, 
         nx30874, nx30877, nx30880, nx30890, nx30893, nx30895, nx30898, nx30900, 
         nx30902, nx30907, nx30909, nx30912, nx30915, nx30925, nx30928, nx30930, 
         nx30933, nx30935, nx30937, nx30940, nx30944, nx30947, nx30950, nx30953, 
         nx30956, nx30959, nx30962, nx30966, nx30968, nx30970, nx30972, nx30974, 
         nx30976, nx30978, nx30980, nx30990, nx30992, nx30998, nx31002, nx31051, 
         nx31098, nx31119, nx31124, nx31126, nx31128, nx31131, nx31135, nx31141, 
         nx31143, nx31146, nx31150, nx31156, nx31159, nx31161, nx31164, nx31166, 
         nx31171, nx31173, nx31176, nx31179, nx31187, nx31193, nx31196, nx31198, 
         nx31201, nx31203, nx31205, nx31210, nx31212, nx31215, nx31218, nx31228, 
         nx31231, nx31233, nx31236, nx31238, nx31240, nx31245, nx31247, nx31250, 
         nx31253, nx31263, nx31266, nx31268, nx31271, nx31273, nx31275, nx31280, 
         nx31282, nx31285, nx31288, nx31298, nx31301, nx31303, nx31306, nx31308, 
         nx31310, nx31315, nx31317, nx31320, nx31323, nx31333, nx31336, nx31338, 
         nx31341, nx31343, nx31345, nx31350, nx31352, nx31355, nx31358, nx31368, 
         nx31371, nx31373, nx31376, nx31378, nx31380, nx31383, nx31387, nx31390, 
         nx31393, nx31396, nx31399, nx31402, nx31405, nx31409, nx31411, nx31413, 
         nx31415, nx31417, nx31419, nx31421, nx31423, nx31429, nx31431, nx31437, 
         nx31441, nx31490, nx31537, nx31558, nx31563, nx31565, nx31567, nx31570, 
         nx31574, nx31580, nx31582, nx31585, nx31589, nx31595, nx31598, nx31600, 
         nx31603, nx31605, nx31610, nx31612, nx31615, nx31618, nx31626, nx31632, 
         nx31635, nx31637, nx31640, nx31642, nx31644, nx31649, nx31651, nx31654, 
         nx31657, nx31667, nx31670, nx31672, nx31675, nx31677, nx31679, nx31684, 
         nx31686, nx31689, nx31692, nx31702, nx31705, nx31707, nx31710, nx31712, 
         nx31714, nx31719, nx31721, nx31724, nx31727, nx31737, nx31740, nx31742, 
         nx31745, nx31747, nx31749, nx31754, nx31756, nx31759, nx31762, nx31772, 
         nx31775, nx31777, nx31780, nx31782, nx31784, nx31789, nx31791, nx31794, 
         nx31797, nx31807, nx31810, nx31812, nx31815, nx31817, nx31819, nx31822, 
         nx31826, nx31829, nx31832, nx31835, nx31838, nx31841, nx31844, nx31848, 
         nx31850, nx31852, nx31854, nx31856, nx31858, nx31860, nx31862, nx31867, 
         nx31869, nx31872, nx31882, nx31893, nx31904, nx31915, nx31926, nx31937, 
         nx31948, nx31959, nx31961, nx31964, nx31974, nx31975, nx31979, nx31989, 
         nx31990, nx31994, nx32004, nx32005, nx32009, nx32019, nx32020, nx32024, 
         nx32034, nx32035, nx32039, nx32049, nx32050, nx32054, nx32056, nx32059, 
         nx32061, nx32071, nx32082, nx32093, nx32104, nx32115, nx32126, nx32137, 
         nx32148, nx32150, nx32153, nx32163, nx32164, nx32168, nx32178, nx32179, 
         nx32183, nx32193, nx32194, nx32198, nx32208, nx32209, nx32213, nx32223, 
         nx32224, nx32228, nx32238, nx32239, nx32243, nx32245, nx32248, nx32252, 
         nx32254, nx32256, nx32259, nx32261, nx32263, nx32266, nx32270, nx32272, 
         nx32276, nx32280, nx32282, nx32284, nx32287, nx32289, nx32291, nx32294, 
         nx32298, nx32300, nx32304, nx32308, nx32310, nx32312, nx32315, nx32317, 
         nx32319, nx32322, nx32326, nx32328, nx32332, nx32336, nx32338, nx32340, 
         nx32343, nx32345, nx32347, nx32350, nx32354, nx32356, nx32360, nx32364, 
         nx32366, nx32368, nx32371, nx32373, nx32375, nx32378, nx32382, nx32384, 
         nx32388, nx32392, nx32394, nx32396, nx32399, nx32401, nx32403, nx32406, 
         nx32410, nx32412, nx32418, nx32420, nx32422, nx32425, nx32427, nx32433, 
         nx32435, nx32446, nx32451, nx32453, nx32464, nx32470, nx32472, nx32475, 
         nx32486, nx32497, nx32508, nx32519, nx32530, nx32541, nx32552, nx32563, 
         nx32565, nx32568, nx32578, nx32579, nx32583, nx32593, nx32594, nx32598, 
         nx32608, nx32609, nx32613, nx32623, nx32624, nx32628, nx32638, nx32639, 
         nx32643, nx32653, nx32654, nx32658, nx32660, nx32665, nx32669, nx32671, 
         nx32682, nx32693, nx32704, nx32715, nx32726, nx32737, nx32748, nx32759, 
         nx32761, nx32764, nx32774, nx32775, nx32779, nx32789, nx32790, nx32794, 
         nx32804, nx32805, nx32809, nx32819, nx32820, nx32824, nx32834, nx32835, 
         nx32839, nx32849, nx32850, nx32854, nx32856, nx32861, nx32865, nx32869, 
         nx32871, nx32880, nx32883, nx32892, nx32894, nx32897, nx32904, nx32908, 
         nx32910, nx32917, nx32921, nx32925, nx32927, nx32936, nx32939, nx32948, 
         nx32950, nx32953, nx32960, nx32964, nx32966, nx32973, nx32977, nx32981, 
         nx32983, nx32992, nx32995, nx33004, nx33006, nx33009, nx33016, nx33020, 
         nx33022, nx33029, nx33033, nx33037, nx33039, nx33048, nx33051, nx33060, 
         nx33062, nx33065, nx33072, nx33076, nx33078, nx33085, nx33089, nx33093, 
         nx33095, nx33104, nx33107, nx33116, nx33118, nx33121, nx33128, nx33132, 
         nx33134, nx33141, nx33145, nx33149, nx33151, nx33160, nx33163, nx33172, 
         nx33174, nx33177, nx33184, nx33188, nx33190, nx33197, nx33203, nx33205, 
         nx33214, nx33217, nx33226, nx33232, nx33234, nx33246, nx33257, nx33259, 
         nx33271, nx33288, nx33290, nx33292, nx33305, nx33316, nx33327, nx33338, 
         nx33349, nx33360, nx33371, nx33382, nx33384, nx33387, nx33397, nx33398, 
         nx33402, nx33412, nx33413, nx33417, nx33427, nx33428, nx33432, nx33442, 
         nx33443, nx33447, nx33457, nx33458, nx33462, nx33472, nx33473, nx33477, 
         nx33479, nx33503, nx33514, nx33525, nx33536, nx33547, nx33558, nx33569, 
         nx33580, nx33582, nx33585, nx33595, nx33596, nx33600, nx33610, nx33611, 
         nx33615, nx33625, nx33626, nx33630, nx33640, nx33641, nx33645, nx33655, 
         nx33656, nx33660, nx33670, nx33671, nx33675, nx33677, nx33694, nx33726, 
         nx33729, nx33731, nx33767, nx33799, nx33802, nx33804, nx33840, nx33872, 
         nx33875, nx33877, nx33913, nx33945, nx33948, nx33950, nx33986, nx34018, 
         nx34021, nx34023, nx34059, nx34091, nx34094, nx34096, nx34162, nx34165, 
         nx34182, nx34209, nx34359, nx34365, nx34368, nx34377, nx34380, nx34389, 
         nx34391, nx34393, nx34395, nx34397, nx34399, nx34401, nx34403, nx34405, 
         nx34407, nx34409, nx34419, nx34429, nx34457, nx34459, nx34461, nx34463, 
         nx34465, nx34467, nx34469, nx34471, nx34473, nx34475, nx34477, nx34479, 
         nx34481, nx34483, nx34485, nx34487, nx34489, nx34491, nx34493, nx34495, 
         nx34499, nx34501, nx34503, nx34505, nx34507, nx34509, nx34511, nx34513, 
         nx34515, nx34517, nx34519, nx34521, nx34523, nx34525, nx34527, nx34529, 
         nx34531, nx34533, nx34535, nx34537, nx34539, nx34541, nx34543, nx34545, 
         nx34547, nx34549, nx34551, nx34553, nx34555, nx34557, nx34571, nx34579, 
         nx34581, nx34583, nx34585, nx34587, nx34589, nx34603, nx34611, nx34613, 
         nx34615, nx34617, nx34619, nx34621, nx34635, nx34643, nx34645, nx34647, 
         nx34649, nx34651, nx34653, nx34667, nx34675, nx34677, nx34679, nx34681, 
         nx34683, nx34705, nx34735, nx34737, nx34739, nx34741, nx34743, nx34745, 
         nx34747, nx34749, nx34751, nx34753, nx34755, nx34757, nx34759, nx34761, 
         nx34763, nx34765, nx34767, nx34769, nx34771, nx34773, nx34775, nx34777, 
         nx34779, nx34781, nx34783, nx34785, nx34787, nx34789, nx34791, nx34793, 
         nx34795, nx34797, nx34799, nx34801, nx34803, nx34805, nx34807, nx34809, 
         nx34811, nx34813, nx34815, nx34817, nx34819, nx34821, nx34833, nx34847, 
         nx34855, nx34857, nx34859, nx34861, nx34863, nx34865, nx34879, nx34887, 
         nx34889, nx34891, nx34893, nx34895, nx34905, nx34913, nx34925, nx34939, 
         nx34947, nx34949, nx34951, nx34953, nx34955, nx34957, nx34971, nx34979, 
         nx34981, nx34983, nx34985, nx34987, nx34997, nx35011, nx35019, nx35021, 
         nx35023, nx35025, nx35027, nx35029, nx35043, nx35051, nx35053, nx35055, 
         nx35057, nx35059, nx35095, nx35097, nx35099, nx35101, nx35103, nx35149, 
         nx35153, nx35155, nx35157, nx35159, nx35161, nx35163, nx35165, nx35167, 
         nx35169, nx35171, nx35173, nx35175, nx35177, nx35179, nx35181, nx35183, 
         nx35185, nx35187, nx35189, nx35191, nx35193, nx35195, nx35197, nx35199, 
         nx35201, nx35205, nx35207, nx35209, nx35211, nx35213, nx35215, nx35217, 
         nx35263, nx35265, nx35267, nx35269, nx35271, nx35289, nx35301, nx35303, 
         nx35305, nx35307, nx35309, nx35313, nx35315, nx35317, nx35319, nx35321, 
         nx35323, nx35325, nx35327, nx35329, nx35331, nx35333, nx35335, nx35339, 
         nx35341, nx35343, nx35345, nx35347, nx35349, nx35351, nx35361, nx35363, 
         nx35365, nx35367, nx35369, nx35371, nx35373, nx35375, nx35377, nx35379, 
         nx35381, nx35385, nx35387, nx35389, nx35391, nx35393, nx35395, nx35397, 
         nx35399, nx35401, nx35403, nx35405, nx35407, nx35411, nx35413, nx35415, 
         nx35417, nx35419, nx35421, nx35423, nx35425, nx35427, nx35429, nx35431, 
         nx35433, nx35437, nx35439, nx35441, nx35443, nx35445, nx35447, nx35449, 
         nx35453, nx35455, nx35457, nx35459, nx35461, nx35463, nx35465, nx35467, 
         nx35469, nx35473, nx35475, nx35477, nx35479, nx35481, nx35485, nx35487, 
         nx35489, nx35491, nx35493, nx35495, nx35497, nx35499, nx35501, nx35503, 
         nx35505, nx35507, nx35511, nx35513, nx35515, nx35517, nx35519, nx35521, 
         nx35523, nx35525, nx35527, nx35529, nx35531, nx35533, nx35537, nx35539, 
         nx35541, nx35543, nx35545, nx35547, nx35549, nx35551, nx35553, nx35555, 
         nx35557, nx35559, nx35563, nx35565, nx35567, nx35569, nx35571, nx35573, 
         nx35575, nx35589, nx35591, nx35593, nx35595, nx35597, nx35599, nx35601, 
         nx35603, nx35605, nx35607, nx35609, nx35615, nx35621, nx35623, nx35625, 
         nx35627, nx35629, nx35631, nx35633, nx35635, nx35637, nx35639, nx35641, 
         nx35643, nx35645, nx35647, nx35649, nx35651, nx35653, nx35655, nx35657, 
         nx35659, nx35661, nx35663, nx35665, nx35667, nx35669, nx35671, nx35673, 
         nx35675, nx35677, nx35679, nx35681, nx35683, nx35685, nx35687, nx35689, 
         nx35691, nx35693, nx35695, nx35697, nx35699, nx35701, nx35703, nx35705, 
         nx35707, nx35709, nx35711, nx35713, nx35715, nx35717, nx35719, nx35721, 
         nx35723, nx35725, nx35727, nx35729, nx35731, nx35733, nx35735, nx35737, 
         nx35739, nx35741, nx35743, nx35745, nx35747, nx35749, nx35751, nx35753, 
         nx35755, nx35757, nx35759, nx35761, nx35763, nx35765, nx35767, nx35769, 
         nx35771, nx35773, nx35775, nx35777, nx35779, nx35781, nx35783, nx35785, 
         nx35787, nx35789, nx35791, nx35793, nx35795, nx35797, nx35799, nx35801, 
         nx35803, nx35805, nx35807, nx35809, nx35811, nx35813, nx35815, nx35817, 
         nx35819, nx35821, nx35823, nx35825, nx35827, nx35829, nx35831, nx35833, 
         nx35835, nx35837, nx35839, nx35841, nx35843, nx35845, nx35847, nx35849, 
         nx35851, nx35853, nx35855, nx35857, nx35859, nx35861, nx35863, nx35865, 
         nx35867, nx35869, nx35871, nx35873, nx35875, nx35877, nx35879, nx35881, 
         nx35883, nx35885, nx35887, nx35889, nx35891, nx35893, nx35895, nx35897, 
         nx35899, nx35901, nx35903, nx35905, nx35907, nx35909, nx35911, nx35913, 
         nx35915, nx35917, nx35919, nx35921, nx35923, nx35925, nx35927, nx35929, 
         nx35931, nx35933, nx35935, nx35937, nx35939, nx35941, nx35943, nx35945, 
         nx35947, nx35949, nx35951, nx35953, nx35955, nx35957, nx35959, nx35961, 
         nx35963, nx35965, nx35967, nx35969, nx35971, nx35973, nx35975, nx35977, 
         nx35979, nx35981, nx35983, nx35985, nx35987, nx35989, nx35991, nx35993, 
         nx35995, nx35997, nx35999, nx36001, nx36003, nx36005, nx36007, nx36009, 
         nx36011, nx36013, nx36015, nx36017, nx36019, nx36021, nx36023, nx36025, 
         nx36027, nx36029, nx36031, nx36033, nx36035, nx36037, nx36039, nx36041, 
         nx36043, nx36045, nx36047, nx36049, nx36051, nx36053, nx36055, nx36057, 
         nx36059, nx36061, nx36063, nx36065, nx36067, nx36069, nx36071, nx36073, 
         nx36075, nx36077, nx36079, nx36081, nx36083, nx36085, nx36087, nx36089, 
         nx36091, nx36093, nx36095, nx36097, nx36099, nx36101, nx36103, nx36105, 
         nx36107, nx36109, nx36111, nx36113, nx36115, nx36117, nx36119, nx36121, 
         nx36123, nx36125, nx36127, nx36129, nx36131, nx36133, nx36135, nx36137, 
         nx36139, nx36141, nx36143, nx36145, nx36147, nx36149, nx36151, nx36153, 
         nx36155, nx36157, nx36159, nx36161, nx36163, nx36165, nx36167, nx36169, 
         nx36171, nx36173, nx36175, nx36177, nx36179, nx36181, nx36183, nx36185, 
         nx36187, nx36189, nx36191, nx36193, nx36195, nx36197, nx36199, nx36201, 
         nx36203, nx36205, nx36207, nx36209, nx36211, nx36213, nx36215, nx36217, 
         nx36219, nx36221, nx36223, nx36225, nx36227, nx36229, nx36231, nx36233, 
         nx36235, nx36237, nx36239, nx36241, nx36243, nx36245, nx36247, nx36249, 
         nx36251, nx36253, nx36255, nx36257, nx36259, nx36261, nx36263, nx36265, 
         nx36267, nx36269, nx36271, nx36273, nx36275, nx36277, nx36279, nx36281, 
         nx36283, nx36285, nx36287, nx36289, nx36291, nx36293, nx36295, nx36297, 
         nx36299, nx36301, nx36307, nx36309, nx36311, nx36313, nx36315, nx36317, 
         nx36319, nx36321, nx36323, nx36325, nx36327, nx36329, nx36331, nx36333, 
         nx36335, nx36337, nx36339, nx36341, nx36343, nx36345, nx36347, nx36349, 
         nx36351, nx36353, nx36355, nx36357, nx36359, nx36361, nx36363, nx36365, 
         nx36367, nx36369, nx36371, nx36373, nx36375, nx36377, nx36379, nx36381, 
         nx36383, nx36385, nx36387, nx36389, nx36391, nx36393;
    wire [800:0] \$dummy ;




    assign enable_write = initiate ;
    fake_vcc ix25758 (.Y (nx25757)) ;
    dffr booth_shift_Reg_adder_0_reg_count_18 (.Q (enable_decoder_dst_booth), .QB (
         \$dummy [0]), .D (nx13613), .CLK (clk), .R (nx34461)) ;
    dffr booth_shift_Reg_adder_0_reg_count_17 (.Q (
         booth_shift_Reg_adder_0_output_17), .QB (\$dummy [1]), .D (nx13603), .CLK (
         clk), .R (nx34461)) ;
    dffr booth_shift_Reg_adder_0_reg_count_16 (.Q (
         booth_shift_Reg_adder_0_output_16), .QB (\$dummy [2]), .D (nx13593), .CLK (
         clk), .R (nx34461)) ;
    dffr booth_shift_Reg_adder_0_reg_count_15 (.Q (
         booth_shift_Reg_adder_0_output_15), .QB (\$dummy [3]), .D (nx13583), .CLK (
         clk), .R (nx34461)) ;
    dffr booth_shift_Reg_adder_0_reg_count_14 (.Q (
         booth_shift_Reg_adder_0_output_14), .QB (\$dummy [4]), .D (nx13573), .CLK (
         clk), .R (nx34461)) ;
    dffr booth_shift_Reg_adder_0_reg_count_13 (.Q (
         booth_shift_Reg_adder_0_output_13), .QB (\$dummy [5]), .D (nx13563), .CLK (
         clk), .R (nx34461)) ;
    dffr booth_shift_Reg_adder_0_reg_count_12 (.Q (
         booth_shift_Reg_adder_0_output_12), .QB (\$dummy [6]), .D (nx13553), .CLK (
         clk), .R (nx34459)) ;
    dffr booth_shift_Reg_adder_0_reg_count_11 (.Q (
         booth_shift_Reg_adder_0_output_11), .QB (\$dummy [7]), .D (nx13543), .CLK (
         clk), .R (nx34459)) ;
    dffr booth_shift_Reg_adder_0_reg_count_10 (.Q (
         booth_shift_Reg_adder_0_output_10), .QB (\$dummy [8]), .D (nx13533), .CLK (
         clk), .R (nx34459)) ;
    dffr booth_shift_Reg_adder_0_reg_count_9 (.Q (
         booth_shift_Reg_adder_0_output_9), .QB (\$dummy [9]), .D (nx13523), .CLK (
         clk), .R (nx34459)) ;
    dffr booth_shift_Reg_adder_0_reg_count_8 (.Q (
         booth_shift_Reg_adder_0_output_8), .QB (\$dummy [10]), .D (nx13513), .CLK (
         clk), .R (nx34459)) ;
    dffr booth_shift_Reg_adder_0_reg_count_7 (.Q (
         booth_shift_Reg_adder_0_output_7), .QB (\$dummy [11]), .D (nx13503), .CLK (
         clk), .R (nx34459)) ;
    dffr booth_shift_Reg_adder_0_reg_count_6 (.Q (
         booth_shift_Reg_adder_0_output_6), .QB (\$dummy [12]), .D (nx13493), .CLK (
         clk), .R (nx34459)) ;
    dffr booth_shift_Reg_adder_0_reg_count_5 (.Q (
         booth_shift_Reg_adder_0_output_5), .QB (\$dummy [13]), .D (nx13483), .CLK (
         clk), .R (nx35615)) ;
    dffr booth_shift_Reg_adder_0_reg_count_4 (.Q (
         booth_shift_Reg_adder_0_output_4), .QB (\$dummy [14]), .D (nx13473), .CLK (
         clk), .R (nx35615)) ;
    dffr booth_shift_Reg_adder_0_reg_count_3 (.Q (
         booth_shift_Reg_adder_0_output_3), .QB (\$dummy [15]), .D (nx13463), .CLK (
         clk), .R (nx35615)) ;
    dffr booth_shift_Reg_adder_0_reg_count_2 (.Q (
         booth_shift_Reg_adder_0_output_2), .QB (\$dummy [16]), .D (nx13453), .CLK (
         clk), .R (nx35615)) ;
    dffr booth_shift_Reg_adder_0_reg_count_1 (.Q (
         booth_shift_Reg_adder_0_output_1), .QB (\$dummy [17]), .D (nx13443), .CLK (
         clk), .R (nx35615)) ;
    dffs_ni booth_shift_Reg_adder_0_reg_count_0 (.Q (
            booth_shift_Reg_adder_0_output_0), .QB (\$dummy [18]), .D (nx13429)
            , .CLK (clk), .S (nx35615)) ;
    dffr reg_ready_signal (.Q (ready_signal), .QB (\$dummy [19]), .D (nx13423), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix14104 (.Y (nx14103), .A0 (state[0]), .A1 (nx830), .S0 (nx12877)
             ) ;
    nor03_2x ix517 (.Y (nx516), .A0 (num_out_2), .A1 (num_out_0), .A2 (num_out_1
             )) ;
    dffr num_loop1_2_fx_reg_q (.Q (num_out_2), .QB (\$dummy [20]), .D (nx13833)
         , .CLK (clk), .R (rst)) ;
    dff reg_num_in_2 (.Q (num_in_2), .QB (\$dummy [21]), .D (nx13823), .CLK (clk
        )) ;
    mux21_ni ix13824 (.Y (nx13823), .A0 (nx496), .A1 (num_in_2), .S0 (nx35161)
             ) ;
    xnor2 ix25822 (.Y (nx25821), .A0 (nx25823), .A1 (nx25986)) ;
    aoi22 ix25824 (.Y (nx25823), .A0 (nx34501), .A1 (alu_inp1_1), .B0 (nx412), .B1 (
          nx12898)) ;
    nand03 ix25828 (.Y (nx25827), .A0 (nx278), .A1 (nx25940), .A2 (nx26129)) ;
    nand02 ix279 (.Y (nx278), .A0 (nx25830), .A1 (nx12887)) ;
    aoi32 ix25831 (.Y (nx25830), .A0 (nx25832), .A1 (nx12882), .A2 (nx266), .B0 (
          nx25900), .B1 (nx258)) ;
    nand02 ix25833 (.Y (nx25832), .A0 (nx12891), .A1 (nx12879)) ;
    nor04_2x ix789 (.Y (nx12891), .A0 (nx25835), .A1 (num_out_3), .A2 (num_out_4
             ), .A3 (nx26044)) ;
    dffr num_loop1_0_fx_reg_q (.Q (num_out_0), .QB (\$dummy [22]), .D (nx13713)
         , .CLK (clk), .R (rst)) ;
    dff reg_num_in_0 (.Q (num_in_0), .QB (\$dummy [23]), .D (nx13703), .CLK (clk
        )) ;
    mux21_ni ix13704 (.Y (nx13703), .A0 (nx376), .A1 (num_in_0), .S0 (nx35159)
             ) ;
    mux21_ni ix13644 (.Y (nx13643), .A0 (nx34393), .A1 (nx210), .S0 (nx12877)) ;
    nand03 ix211 (.Y (nx210), .A0 (nx25849), .A1 (nx35103), .A2 (nx35149)) ;
    nand02 ix25850 (.Y (nx25849), .A0 (nx25813), .A1 (nx12879)) ;
    dffr reg_state_1 (.Q (state[1]), .QB (\$dummy [24]), .D (nx13643), .CLK (clk
         ), .R (rst)) ;
    nand02 ix25855 (.Y (nx25854), .A0 (nx34397), .A1 (nx172)) ;
    dffr reg_state_0 (.Q (state[0]), .QB (nx25857), .D (nx14103), .CLK (clk), .R (
         rst)) ;
    dffr reg_state_2 (.Q (state[2]), .QB (\$dummy [25]), .D (nx14093), .CLK (clk
         ), .R (rst)) ;
    dff reg_alu_inp1_0 (.Q (alu_inp1_0), .QB (\$dummy [26]), .D (nx13723), .CLK (
        clk)) ;
    mux21_ni ix13724 (.Y (nx13723), .A0 (nx390), .A1 (alu_inp1_0), .S0 (nx35095)
             ) ;
    dffr address_loop1_0_fx_reg_q (.Q (address_out_0), .QB (\$dummy [27]), .D (
         nx13693), .CLK (clk), .R (rst)) ;
    mux21_ni ix13694 (.Y (nx13693), .A0 (address_out_0), .A1 (address_in_0), .S0 (
             nx34503)) ;
    dffr reg_address_in_0 (.Q (address_in_0), .QB (\$dummy [28]), .D (nx13683), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix13684 (.Y (nx13683), .A0 (address_in_0), .A1 (nx358), .S0 (
             nx34507)) ;
    nor02_2x ix359 (.Y (nx358), .A0 (nx25864), .A1 (nx35787)) ;
    dffr reg_sub_state_1 (.Q (sub_state[1]), .QB (\$dummy [29]), .D (nx13413), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix13414 (.Y (nx13413), .A0 (sub_state[1]), .A1 (nx26), .S0 (nx12883
             )) ;
    oai21 ix25880 (.Y (nx25879), .A0 (sub_state[1]), .A1 (nx34401), .B0 (nx35157
          )) ;
    dffr reg_sub_state_0 (.Q (sub_state[0]), .QB (\$dummy [30]), .D (nx13403), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix13404 (.Y (nx13403), .A0 (nx34401), .A1 (nx20), .S0 (nx12883)) ;
    oai22 ix183 (.Y (nx12883), .A0 (nx35155), .A1 (nx25891), .B0 (nx12879), .B1 (
          nx25893)) ;
    nand02 ix25892 (.Y (nx25891), .A0 (nx25813), .A1 (nx12879)) ;
    aoi21 ix25897 (.Y (nx25896), .A0 (sub_state[1]), .A1 (nx34401), .B0 (nx34397
          )) ;
    oai43 ix351 (.Y (nx350), .A0 (nx35155), .A1 (nx12891), .A2 (nx25900), .A3 (
          nx25902), .B0 (nx25919), .B1 (nx34389), .B2 (nx34393)) ;
    oai21 ix25903 (.Y (nx25902), .A0 (nx334), .A1 (nx25916), .B0 (nx258)) ;
    nor02_2x ix259 (.Y (nx258), .A0 (nx34401), .A1 (nx25879)) ;
    dffr reg_sub_state_2 (.Q (sub_state[2]), .QB (\$dummy [31]), .D (nx13633), .CLK (
         clk), .R (rst)) ;
    xnor2 ix321 (.Y (nx320), .A0 (sub_state[1]), .A1 (nx34401)) ;
    dff reg_enable_address (.Q (enable_address), .QB (\$dummy [32]), .D (nx13673
        ), .CLK (clk)) ;
    or02 ix13674 (.Y (nx13673), .A0 (nx34503), .A1 (nx300)) ;
    nor03_2x ix301 (.Y (nx300), .A0 (nx38), .A1 (rst), .A2 (nx35099)) ;
    nand02 ix39 (.Y (nx38), .A0 (nx35157), .A1 (nx34401)) ;
    nand02 ix13734 (.Y (nx13733), .A0 (nx25935), .A1 (nx35095)) ;
    dff reg_alu_inp2_0 (.Q (\$dummy [33]), .QB (nx25935), .D (nx13733), .CLK (
        clk)) ;
    nand03 ix25938 (.Y (nx25937), .A0 (nx242), .A1 (nx25940), .A2 (nx25942)) ;
    inv01 ix25941 (.Y (nx25940), .A (rst)) ;
    nand02 ix25943 (.Y (nx25942), .A0 (nx25944), .A1 (nx34405)) ;
    nor03_2x ix25945 (.Y (nx25944), .A0 (sub_state[1]), .A1 (nx34403), .A2 (
             nx34397)) ;
    nand02 ix13654 (.Y (nx13653), .A0 (nx35795), .A1 (nx25951)) ;
    dffr reg_enable_num (.Q (\$dummy [34]), .QB (nx25949), .D (nx13653), .CLK (
         clk), .R (rst)) ;
    nand02 ix25952 (.Y (nx25951), .A0 (nx34495), .A1 (nx25944)) ;
    dffr num_loop1_1_fx_reg_q (.Q (num_out_1), .QB (\$dummy [35]), .D (nx13773)
         , .CLK (clk), .R (rst)) ;
    mux21 ix13764 (.Y (nx13763), .A0 (nx25958), .A1 (nx25975), .S0 (nx35159)) ;
    aoi22 ix25959 (.Y (nx25958), .A0 (mdr_data_out[1]), .A1 (nx34495), .B0 (
          nx414), .B1 (nx34405)) ;
    xnor2 ix415 (.Y (nx414), .A0 (nx412), .A1 (nx25962)) ;
    dff reg_alu_inp1_1 (.Q (alu_inp1_1), .QB (\$dummy [36]), .D (nx13783), .CLK (
        clk)) ;
    mux21_ni ix13784 (.Y (nx13783), .A0 (nx448), .A1 (alu_inp1_1), .S0 (nx35095)
             ) ;
    dffr address_loop1_1_fx_reg_q (.Q (address_out_1), .QB (\$dummy [37]), .D (
         nx13753), .CLK (clk), .R (rst)) ;
    mux21_ni ix13754 (.Y (nx13753), .A0 (address_out_1), .A1 (address_in_1), .S0 (
             nx34503)) ;
    dffr reg_address_in_1 (.Q (address_in_1), .QB (\$dummy [38]), .D (nx13743), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix13744 (.Y (nx13743), .A0 (address_in_1), .A1 (nx416), .S0 (
             nx34507)) ;
    nor02ii ix417 (.Y (nx416), .A0 (nx35787), .A1 (nx414)) ;
    dff reg_num_in_1 (.Q (num_in_1), .QB (nx25975), .D (nx13763), .CLK (clk)) ;
    dffr num_loop1_3_fx_reg_q (.Q (num_out_3), .QB (\$dummy [39]), .D (nx13883)
         , .CLK (clk), .R (rst)) ;
    mux21 ix13874 (.Y (nx13873), .A0 (nx25982), .A1 (nx26014), .S0 (nx35159)) ;
    aoi22 ix25983 (.Y (nx25982), .A0 (mdr_data_out[3]), .A1 (nx34495), .B0 (
          nx12901), .B1 (nx34405)) ;
    xnor2 ix551 (.Y (nx12901), .A0 (nx522), .A1 (nx26001)) ;
    oai22 ix523 (.Y (nx522), .A0 (nx25823), .A1 (nx25986), .B0 (nx35799), .B1 (
          nx25998)) ;
    dff reg_alu_inp1_2 (.Q (alu_inp1_2), .QB (nx25998), .D (nx13813), .CLK (clk)
        ) ;
    mux21_ni ix13814 (.Y (nx13813), .A0 (nx480), .A1 (alu_inp1_2), .S0 (nx35095)
             ) ;
    dffr address_loop1_2_fx_reg_q (.Q (address_out_2), .QB (\$dummy [40]), .D (
         nx13803), .CLK (clk), .R (rst)) ;
    mux21_ni ix13804 (.Y (nx13803), .A0 (address_out_2), .A1 (address_in_2), .S0 (
             nx34503)) ;
    dffr reg_address_in_2 (.Q (address_in_2), .QB (\$dummy [41]), .D (nx13793), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix13794 (.Y (nx13793), .A0 (address_in_2), .A1 (nx464), .S0 (
             nx34507)) ;
    nor02_2x ix465 (.Y (nx464), .A0 (nx25821), .A1 (nx35787)) ;
    dff reg_alu_sel (.Q (\$dummy [42]), .QB (nx25999), .D (nx13663), .CLK (clk)
        ) ;
    dff reg_alu_inp1_3 (.Q (alu_inp1_3), .QB (\$dummy [43]), .D (nx13863), .CLK (
        clk)) ;
    mux21_ni ix13864 (.Y (nx13863), .A0 (nx540), .A1 (alu_inp1_3), .S0 (nx35095)
             ) ;
    dffr address_loop1_3_fx_reg_q (.Q (address_out_3), .QB (\$dummy [44]), .D (
         nx13853), .CLK (clk), .R (rst)) ;
    mux21_ni ix13854 (.Y (nx13853), .A0 (address_out_3), .A1 (address_in_3), .S0 (
             nx34503)) ;
    dffr reg_address_in_3 (.Q (address_in_3), .QB (\$dummy [45]), .D (nx13843), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix13844 (.Y (nx13843), .A0 (address_in_3), .A1 (nx524), .S0 (
             nx34507)) ;
    nor02ii ix525 (.Y (nx524), .A0 (nx35787), .A1 (nx12901)) ;
    dff reg_num_in_3 (.Q (num_in_3), .QB (nx26014), .D (nx13873), .CLK (clk)) ;
    dffr num_loop1_4_fx_reg_q (.Q (num_out_4), .QB (\$dummy [46]), .D (nx13933)
         , .CLK (clk), .R (rst)) ;
    dff reg_num_in_4 (.Q (num_in_4), .QB (\$dummy [47]), .D (nx13923), .CLK (clk
        )) ;
    mux21_ni ix13924 (.Y (nx13923), .A0 (nx606), .A1 (num_in_4), .S0 (nx35159)
             ) ;
    xnor2 ix26023 (.Y (nx26022), .A0 (nx26024), .A1 (nx26027)) ;
    aoi22 ix26025 (.Y (nx26024), .A0 (nx34499), .A1 (alu_inp1_3), .B0 (nx522), .B1 (
          nx548)) ;
    dff reg_alu_inp1_4 (.Q (alu_inp1_4), .QB (nx26039), .D (nx13913), .CLK (clk)
        ) ;
    mux21_ni ix13914 (.Y (nx13913), .A0 (nx590), .A1 (alu_inp1_4), .S0 (nx35095)
             ) ;
    dffr address_loop1_4_fx_reg_q (.Q (address_out_4), .QB (\$dummy [48]), .D (
         nx13903), .CLK (clk), .R (rst)) ;
    mux21_ni ix13904 (.Y (nx13903), .A0 (address_out_4), .A1 (address_in_4), .S0 (
             nx34503)) ;
    dffr reg_address_in_4 (.Q (address_in_4), .QB (\$dummy [49]), .D (nx13893), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix13894 (.Y (nx13893), .A0 (address_in_4), .A1 (nx574), .S0 (
             nx34507)) ;
    nor02_2x ix575 (.Y (nx574), .A0 (nx26022), .A1 (nx35787)) ;
    dffr num_loop1_5_fx_reg_q (.Q (num_out_5), .QB (nx26046), .D (nx13983), .CLK (
         clk), .R (rst)) ;
    mux21 ix13974 (.Y (nx13973), .A0 (nx26052), .A1 (nx26069), .S0 (nx35159)) ;
    aoi22 ix26053 (.Y (nx26052), .A0 (mdr_data_out[5]), .A1 (nx34495), .B0 (
          nx12905), .B1 (nx34405)) ;
    xnor2 ix659 (.Y (nx12905), .A0 (nx630), .A1 (nx26056)) ;
    oai22 ix631 (.Y (nx630), .A0 (nx26024), .A1 (nx26027), .B0 (nx35799), .B1 (
          nx26039)) ;
    dff reg_alu_inp1_5 (.Q (alu_inp1_5), .QB (\$dummy [50]), .D (nx13963), .CLK (
        clk)) ;
    mux21_ni ix13964 (.Y (nx13963), .A0 (nx648), .A1 (alu_inp1_5), .S0 (nx35095)
             ) ;
    dffr address_loop1_5_fx_reg_q (.Q (address_out_5), .QB (\$dummy [51]), .D (
         nx13953), .CLK (clk), .R (rst)) ;
    mux21_ni ix13954 (.Y (nx13953), .A0 (address_out_5), .A1 (address_in_5), .S0 (
             nx34503)) ;
    dffr reg_address_in_5 (.Q (address_in_5), .QB (\$dummy [52]), .D (nx13943), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix13944 (.Y (nx13943), .A0 (address_in_5), .A1 (nx632), .S0 (
             nx34507)) ;
    nor02ii ix633 (.Y (nx632), .A0 (nx35787), .A1 (nx12905)) ;
    dff reg_num_in_5 (.Q (\$dummy [53]), .QB (nx26069), .D (nx13973), .CLK (clk)
        ) ;
    dffr num_loop1_6_fx_reg_q (.Q (num_out_6), .QB (\$dummy [54]), .D (nx14033)
         , .CLK (clk), .R (rst)) ;
    dff reg_num_in_6 (.Q (num_in_6), .QB (\$dummy [55]), .D (nx14023), .CLK (clk
        )) ;
    mux21_ni ix14024 (.Y (nx14023), .A0 (nx714), .A1 (num_in_6), .S0 (nx35159)
             ) ;
    xnor2 ix26079 (.Y (nx26078), .A0 (nx26080), .A1 (nx26083)) ;
    aoi22 ix26081 (.Y (nx26080), .A0 (nx34501), .A1 (alu_inp1_5), .B0 (nx630), .B1 (
          nx656)) ;
    dff reg_alu_inp1_6 (.Q (alu_inp1_6), .QB (nx26095), .D (nx14013), .CLK (clk)
        ) ;
    mux21_ni ix14014 (.Y (nx14013), .A0 (nx698), .A1 (alu_inp1_6), .S0 (nx35097)
             ) ;
    dffr address_loop1_6_fx_reg_q (.Q (address_out_6), .QB (\$dummy [56]), .D (
         nx14003), .CLK (clk), .R (rst)) ;
    mux21_ni ix14004 (.Y (nx14003), .A0 (address_out_6), .A1 (address_in_6), .S0 (
             nx34505)) ;
    dffr reg_address_in_6 (.Q (address_in_6), .QB (\$dummy [57]), .D (nx13993), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix13994 (.Y (nx13993), .A0 (address_in_6), .A1 (nx682), .S0 (
             nx34507)) ;
    nor02_2x ix683 (.Y (nx682), .A0 (nx26078), .A1 (nx35787)) ;
    dffr num_loop1_7_fx_reg_q (.Q (num_out_7), .QB (nx26099), .D (nx14083), .CLK (
         clk), .R (rst)) ;
    mux21 ix14074 (.Y (nx14073), .A0 (nx26105), .A1 (nx26122), .S0 (nx35159)) ;
    aoi22 ix26106 (.Y (nx26105), .A0 (mdr_data_out[7]), .A1 (nx34495), .B0 (
          nx12907), .B1 (nx34407)) ;
    xnor2 ix765 (.Y (nx12907), .A0 (nx736), .A1 (nx26109)) ;
    oai22 ix737 (.Y (nx736), .A0 (nx26080), .A1 (nx26083), .B0 (nx35799), .B1 (
          nx26095)) ;
    dff reg_alu_inp1_7 (.Q (alu_inp1_7), .QB (\$dummy [58]), .D (nx14063), .CLK (
        clk)) ;
    mux21_ni ix14064 (.Y (nx14063), .A0 (nx754), .A1 (alu_inp1_7), .S0 (nx35097)
             ) ;
    dffr address_loop1_7_fx_reg_q (.Q (address_out_7), .QB (\$dummy [59]), .D (
         nx14053), .CLK (clk), .R (rst)) ;
    mux21_ni ix14054 (.Y (nx14053), .A0 (address_out_7), .A1 (address_in_7), .S0 (
             nx34505)) ;
    dffr reg_address_in_7 (.Q (address_in_7), .QB (\$dummy [60]), .D (nx14043), 
         .CLK (clk), .R (rst)) ;
    mux21_ni ix14044 (.Y (nx14043), .A0 (address_in_7), .A1 (nx738), .S0 (
             nx34509)) ;
    nor02ii ix739 (.Y (nx738), .A0 (nx35789), .A1 (nx12907)) ;
    dff reg_num_in_7 (.Q (\$dummy [61]), .QB (nx26122), .D (nx14073), .CLK (clk)
        ) ;
    dffr booth_shift_Reg_adder_0_reg_count_19 (.Q (done), .QB (\$dummy [62]), .D (
         nx13623), .CLK (clk), .R (nx35615)) ;
    aoi21 ix267 (.Y (nx266), .A0 (nx34403), .A1 (nx174), .B0 (nx38)) ;
    aoi21 ix807 (.Y (nx12887), .A0 (nx34395), .A1 (state[0]), .B0 (nx34391)) ;
    aoi21 ix26130 (.Y (nx26129), .A0 (nx25942), .A1 (nx846), .B0 (nx12909)) ;
    nand02 ix57 (.Y (nx56), .A0 (nx26144), .A1 (nx25832)) ;
    oai21 ix26145 (.Y (nx26144), .A0 (nx12885), .A1 (nx35155), .B0 (nx12879)) ;
    fake_gnd ix12510 (.Y (initiate)) ;
    dffr max_calc_reg_done_comp (.Q (done_comp), .QB (\$dummy [63]), .D (nx25723
         ), .CLK (clk), .R (rst)) ;
    or02 ix25724 (.Y (nx25723), .A0 (done_comp), .A1 (nx35741)) ;
    oai32 ix17574 (.Y (nx17573), .A0 (nx36389), .A1 (start_comp), .A2 (
          max_calc_start), .B0 (nx26184), .B1 (nx26191)) ;
    dffr max_calc_reg_state_2 (.Q (max_calc_state_2), .QB (\$dummy [64]), .D (
         nx17573), .CLK (clk), .R (rst)) ;
    nand02 ix17524 (.Y (nx17523), .A0 (nx26176), .A1 (nx25832)) ;
    dffr reg_start_comp (.Q (start_comp), .QB (nx26176), .D (nx17523), .CLK (clk
         ), .R (rst)) ;
    nand02 ix17534 (.Y (nx17533), .A0 (nx26180), .A1 (nx26182)) ;
    dffr max_calc_reg_start (.Q (max_calc_start), .QB (nx26180), .D (nx17533), .CLK (
         clk), .R (rst)) ;
    aoi43 ix26185 (.Y (nx26184), .A0 (nx26186), .A1 (nx34705), .A2 (nx36389), .A3 (
          nx26203), .B0 (nx34737), .B1 (nx26182), .B2 (nx26201)) ;
    aoi21 ix26187 (.Y (nx26186), .A0 (nx26188), .A1 (nx6300), .B0 (nx6244)) ;
    dffr max_calc_reg_state_0 (.Q (max_calc_state_0), .QB (nx26188), .D (nx17543
         ), .CLK (clk), .R (rst)) ;
    oai32 ix17544 (.Y (nx17543), .A0 (nx26188), .A1 (start_comp), .A2 (
          max_calc_start), .B0 (nx26186), .B1 (nx26191)) ;
    aoi21 ix6301 (.Y (nx6300), .A0 (nx36389), .A1 (nx26194), .B0 (
          max_calc_state_3)) ;
    dffr max_calc_reg_state_3 (.Q (max_calc_state_3), .QB (nx26203), .D (nx17563
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_state_1 (.Q (max_calc_state_1), .QB (\$dummy [65]), .D (
         nx17553), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_0 (.Q (answer[0]), .QB (\$dummy [66]), .D (nx25563)
         , .CLK (clk), .R (rst)) ;
    dff max_calc_reg_comparator_first_inp1_0 (.Q (
        max_calc_comparator_first_inp1_0), .QB (\$dummy [67]), .D (nx19633), .CLK (
        clk)) ;
    dffr labelsregfile_label1_loop1_0_fx_reg_q (.Q (label_1_output[0]), .QB (
         \$dummy [68]), .D (nx17223), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_0 (.Q (label_1_input_0), .D (nx5758), .CLK (nx34511)
          ) ;
    oai21 ix5759 (.Y (nx5758), .A0 (nx26223), .A1 (nx34409), .B0 (nx26227)) ;
    dffr reg_label_1_input_state_machine_0 (.Q (label_1_input_state_machine_0), 
         .QB (nx26223), .D (nx17213), .CLK (clk), .R (rst)) ;
    oai21 ix26228 (.Y (nx26227), .A0 (nx35731), .A1 (label_1_output[0]), .B0 (
          nx5746)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_0_1), .QB (\$dummy [69]), .D (nx17193), 
         .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_0_2), .QB (nx26648), .D (nx17183), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_0_3), .QB (\$dummy [70]), .D (nx17173), 
         .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_0_4), .QB (nx26646), .D (nx17163), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_0_5), .QB (\$dummy [71]), .D (nx17153), 
         .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_0_6), .QB (nx26644), .D (nx17143), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_0_7), .QB (\$dummy [72]), .D (nx17133), 
         .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_0_8), .QB (nx26642), .D (nx17123), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_0_9), .QB (\$dummy [73]), .D (nx17113), 
         .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_0_10), .QB (nx26640), .D (nx17103), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_0_11), .QB (\$dummy [74]), .D (nx17093)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_0_12), .QB (nx26638), .D (nx17083), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_0_13), .QB (\$dummy [75]), .D (nx17073)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_0_14), .QB (nx26636), .D (nx17063), .CLK (
         clk), .R (rst)) ;
    aoi22 ix26277 (.Y (nx26276), .A0 (mdr_data_out[15]), .A1 (nx34667), .B0 (
          nx5544), .B1 (nx5550)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_reg_output_0), .QB (\$dummy [76]), .D (
         nx16703), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_0_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_0_shift_Reg_count_0), .QB (\$dummy [77]), .D (
            nx16689), .CLK (clk), .S (nx34465)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_reg_output_9), .QB (\$dummy [78]), .D (
         nx16883), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_9), .QB (\$dummy [79]), .D (
         nx16873), .CLK (clk), .R (nx34465)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_8), .QB (\$dummy [80]), .D (
         nx16863), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_8), .QB (\$dummy [81]), .D (
         nx16853), .CLK (clk), .R (nx34465)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_7), .QB (\$dummy [82]), .D (
         nx16843), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_7), .QB (\$dummy [83]), .D (
         nx16833), .CLK (clk), .R (nx34463)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_6), .QB (\$dummy [84]), .D (
         nx16823), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_6), .QB (\$dummy [85]), .D (
         nx16813), .CLK (clk), .R (nx34463)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_5), .QB (\$dummy [86]), .D (
         nx16803), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_5), .QB (\$dummy [87]), .D (
         nx16793), .CLK (clk), .R (nx34463)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_4), .QB (\$dummy [88]), .D (
         nx16783), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_4), .QB (\$dummy [89]), .D (
         nx16773), .CLK (clk), .R (nx34463)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_3), .QB (\$dummy [90]), .D (
         nx16763), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_3), .QB (\$dummy [91]), .D (
         nx16753), .CLK (clk), .R (nx34463)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_2), .QB (\$dummy [92]), .D (
         nx16743), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_2), .QB (\$dummy [93]), .D (
         nx16733), .CLK (clk), .R (nx34463)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_0_shift_Reg_output_1), .QB (\$dummy [94]), .D (
         nx16723), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_0_shift_Reg_count_1), .QB (\$dummy [95]), .D (
         nx16713), .CLK (clk), .R (nx34461)) ;
    nand02 ix16684 (.Y (nx16683), .A0 (nx35803), .A1 (nx34653)) ;
    dffs_ni booth_booth_integrtaion_0_shift_Reg_reg_en (.Q (\$dummy [96]), .QB (
            nx26323), .D (nx16683), .CLK (clk), .S (nx34463)) ;
    nand02 ix5545 (.Y (nx5544), .A0 (nx26344), .A1 (nx26356)) ;
    oai21 ix26345 (.Y (nx26344), .A0 (nx34681), .A1 (nx34675), .B0 (
          mdr_data_out[16])) ;
    oai21 ix16894 (.Y (nx16893), .A0 (nx26349), .A1 (nx35193), .B0 (nx26351)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [97]), .QB (
         nx26349), .D (nx16893), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [98]), .QB (
         nx26353), .D (nx17203), .CLK (clk), .R (rst)) ;
    xnor2 ix26361 (.Y (nx26360), .A0 (nx5014), .A1 (nx13067)) ;
    oai21 ix17034 (.Y (nx17033), .A0 (nx26366), .A1 (nx35193), .B0 (nx26368)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_17), .QB (nx26366), .D (nx17033)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26369 (.Y (nx26368), .A0 (nx35201), .A1 (nx5522), .A2 (nx36003)) ;
    xnor2 ix5523 (.Y (nx5522), .A0 (nx26371), .A1 (nx13069)) ;
    aoi22 ix26372 (.Y (nx26371), .A0 (booth_booth_integrtaion_0_booth_output_17)
          , .A1 (nx5038), .B0 (nx5014), .B1 (nx13067)) ;
    nand02 ix5023 (.Y (nx5022), .A0 (mdr_data_out[17]), .A1 (mdr_data_out[16])
           ) ;
    or02 ix26376 (.Y (nx26375), .A0 (mdr_data_out[16]), .A1 (mdr_data_out[17])
         ) ;
    xnor2 ix26382 (.Y (nx26381), .A0 (nx5066), .A1 (nx13071)) ;
    oai22 ix5067 (.Y (nx5066), .A0 (nx26371), .A1 (nx26384), .B0 (nx26391), .B1 (
          nx35205)) ;
    aoi32 ix26387 (.Y (nx26386), .A0 (nx5048), .A1 (nx34681), .A2 (nx26389), .B0 (
          mdr_data_out[18]), .B1 (nx34675)) ;
    oai21 ix5049 (.Y (nx5048), .A0 (mdr_data_out[16]), .A1 (mdr_data_out[17]), .B0 (
          mdr_data_out[18])) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_18), .QB (nx26391), .D (nx17023)
         , .CLK (clk), .R (rst)) ;
    oai21 ix17014 (.Y (nx17013), .A0 (nx26396), .A1 (nx35193), .B0 (nx26398)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_19), .QB (nx26396), .D (nx17013)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26399 (.Y (nx26398), .A0 (nx35201), .A1 (nx5498), .A2 (nx36003)) ;
    xnor2 ix5499 (.Y (nx5498), .A0 (nx26401), .A1 (nx13073)) ;
    aoi22 ix26402 (.Y (nx26401), .A0 (booth_booth_integrtaion_0_booth_output_19)
          , .A1 (nx5086), .B0 (nx5066), .B1 (nx13071)) ;
    nor02ii ix26405 (.Y (nx26404), .A0 (nx5052), .A1 (mdr_data_out[19])) ;
    nor03_2x ix5053 (.Y (nx5052), .A0 (mdr_data_out[18]), .A1 (mdr_data_out[16])
             , .A2 (mdr_data_out[17])) ;
    nor04 ix5077 (.Y (nx5076), .A0 (mdr_data_out[19]), .A1 (mdr_data_out[18]), .A2 (
          mdr_data_out[16]), .A3 (mdr_data_out[17])) ;
    xnor2 ix26419 (.Y (nx26418), .A0 (nx5114), .A1 (nx13074)) ;
    oai22 ix5115 (.Y (nx5114), .A0 (nx26401), .A1 (nx26421), .B0 (nx26430), .B1 (
          nx35207)) ;
    aoi32 ix26424 (.Y (nx26423), .A0 (nx5096), .A1 (nx34681), .A2 (nx26428), .B0 (
          mdr_data_out[20]), .B1 (nx34675)) ;
    nand02 ix5097 (.Y (nx5096), .A0 (nx26426), .A1 (mdr_data_out[20])) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_20), .QB (nx26430), .D (nx17003)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16994 (.Y (nx16993), .A0 (nx26435), .A1 (nx35193), .B0 (nx26437)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_21), .QB (nx26435), .D (nx16993)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26438 (.Y (nx26437), .A0 (nx35201), .A1 (nx5474), .A2 (nx36003)) ;
    xnor2 ix5475 (.Y (nx5474), .A0 (nx26440), .A1 (nx13075)) ;
    aoi22 ix26441 (.Y (nx26440), .A0 (booth_booth_integrtaion_0_booth_output_21)
          , .A1 (nx5134), .B0 (nx5114), .B1 (nx13074)) ;
    nor02ii ix26444 (.Y (nx26443), .A0 (nx5100), .A1 (mdr_data_out[21])) ;
    nor02ii ix5101 (.Y (nx5100), .A0 (mdr_data_out[20]), .A1 (nx5076)) ;
    nor02ii ix5125 (.Y (nx5124), .A0 (mdr_data_out[21]), .A1 (nx5100)) ;
    xnor2 ix26454 (.Y (nx26453), .A0 (nx5162), .A1 (nx13077)) ;
    oai22 ix5163 (.Y (nx5162), .A0 (nx26440), .A1 (nx26456), .B0 (nx26465), .B1 (
          nx35209)) ;
    aoi32 ix26459 (.Y (nx26458), .A0 (nx5144), .A1 (nx34681), .A2 (nx26463), .B0 (
          mdr_data_out[22]), .B1 (nx34675)) ;
    nand02 ix5145 (.Y (nx5144), .A0 (nx26461), .A1 (mdr_data_out[22])) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_22), .QB (nx26465), .D (nx16983)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16974 (.Y (nx16973), .A0 (nx26470), .A1 (nx35193), .B0 (nx26472)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_23), .QB (nx26470), .D (nx16973)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26473 (.Y (nx26472), .A0 (nx35201), .A1 (nx5450), .A2 (nx35195)) ;
    xnor2 ix5451 (.Y (nx5450), .A0 (nx26475), .A1 (nx13079)) ;
    aoi22 ix26476 (.Y (nx26475), .A0 (booth_booth_integrtaion_0_booth_output_23)
          , .A1 (nx5182), .B0 (nx5162), .B1 (nx13077)) ;
    nor02ii ix26479 (.Y (nx26478), .A0 (nx5148), .A1 (mdr_data_out[23])) ;
    nor02ii ix5149 (.Y (nx5148), .A0 (mdr_data_out[22]), .A1 (nx5124)) ;
    nor02ii ix5173 (.Y (nx5172), .A0 (mdr_data_out[23]), .A1 (nx5148)) ;
    xnor2 ix26489 (.Y (nx26488), .A0 (nx5210), .A1 (nx13081)) ;
    oai22 ix5211 (.Y (nx5210), .A0 (nx26475), .A1 (nx26491), .B0 (nx26500), .B1 (
          nx35211)) ;
    aoi32 ix26494 (.Y (nx26493), .A0 (nx5192), .A1 (nx34681), .A2 (nx26498), .B0 (
          mdr_data_out[24]), .B1 (nx34675)) ;
    nand02 ix5193 (.Y (nx5192), .A0 (nx26496), .A1 (mdr_data_out[24])) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_24), .QB (nx26500), .D (nx16963)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16954 (.Y (nx16953), .A0 (nx26505), .A1 (nx35195), .B0 (nx26507)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_25), .QB (nx26505), .D (nx16953)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26508 (.Y (nx26507), .A0 (nx35201), .A1 (nx5426), .A2 (nx35195)) ;
    xnor2 ix5427 (.Y (nx5426), .A0 (nx26510), .A1 (nx13083)) ;
    aoi22 ix26511 (.Y (nx26510), .A0 (booth_booth_integrtaion_0_booth_output_25)
          , .A1 (nx5230), .B0 (nx5210), .B1 (nx13081)) ;
    nor02ii ix26514 (.Y (nx26513), .A0 (nx5196), .A1 (mdr_data_out[25])) ;
    nor02ii ix5197 (.Y (nx5196), .A0 (mdr_data_out[24]), .A1 (nx5172)) ;
    nor02ii ix5221 (.Y (nx5220), .A0 (mdr_data_out[25]), .A1 (nx5196)) ;
    xnor2 ix26524 (.Y (nx26523), .A0 (nx5258), .A1 (nx13085)) ;
    oai22 ix5259 (.Y (nx5258), .A0 (nx26510), .A1 (nx26526), .B0 (nx26535), .B1 (
          nx35213)) ;
    aoi32 ix26529 (.Y (nx26528), .A0 (nx5240), .A1 (nx34681), .A2 (nx26533), .B0 (
          mdr_data_out[26]), .B1 (nx34675)) ;
    nand02 ix5241 (.Y (nx5240), .A0 (nx26531), .A1 (mdr_data_out[26])) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_26), .QB (nx26535), .D (nx16943)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16934 (.Y (nx16933), .A0 (nx26540), .A1 (nx35195), .B0 (nx26542)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_27), .QB (nx26540), .D (nx16933)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26543 (.Y (nx26542), .A0 (nx35201), .A1 (nx5402), .A2 (nx35195)) ;
    xnor2 ix5403 (.Y (nx5402), .A0 (nx26545), .A1 (nx13087)) ;
    aoi22 ix26546 (.Y (nx26545), .A0 (booth_booth_integrtaion_0_booth_output_27)
          , .A1 (nx5278), .B0 (nx5258), .B1 (nx13085)) ;
    nor02ii ix26549 (.Y (nx26548), .A0 (nx5244), .A1 (mdr_data_out[27])) ;
    nor02ii ix5245 (.Y (nx5244), .A0 (mdr_data_out[26]), .A1 (nx5220)) ;
    nor02ii ix5269 (.Y (nx5268), .A0 (mdr_data_out[27]), .A1 (nx5244)) ;
    xnor2 ix26559 (.Y (nx26558), .A0 (nx5306), .A1 (nx13089)) ;
    oai22 ix5307 (.Y (nx5306), .A0 (nx26545), .A1 (nx26561), .B0 (nx26570), .B1 (
          nx35215)) ;
    aoi32 ix26564 (.Y (nx26563), .A0 (nx5288), .A1 (nx34681), .A2 (nx26568), .B0 (
          mdr_data_out[28]), .B1 (nx34675)) ;
    nand02 ix5289 (.Y (nx5288), .A0 (nx26566), .A1 (mdr_data_out[28])) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_28), .QB (nx26570), .D (nx16923)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16914 (.Y (nx16913), .A0 (nx26575), .A1 (nx35195), .B0 (nx26577)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_29), .QB (nx26575), .D (nx16913)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26578 (.Y (nx26577), .A0 (nx36011), .A1 (nx5378), .A2 (nx35195)) ;
    xnor2 ix5379 (.Y (nx5378), .A0 (nx26580), .A1 (nx13090)) ;
    aoi22 ix26581 (.Y (nx26580), .A0 (booth_booth_integrtaion_0_booth_output_29)
          , .A1 (nx5326), .B0 (nx5306), .B1 (nx13089)) ;
    nor02ii ix26584 (.Y (nx26583), .A0 (nx5292), .A1 (mdr_data_out[29])) ;
    nor02ii ix5293 (.Y (nx5292), .A0 (mdr_data_out[28]), .A1 (nx5268)) ;
    nor02ii ix5317 (.Y (nx5316), .A0 (mdr_data_out[29]), .A1 (nx5292)) ;
    xnor2 ix26594 (.Y (nx26593), .A0 (nx5354), .A1 (nx5364)) ;
    oai22 ix5355 (.Y (nx5354), .A0 (nx26580), .A1 (nx26596), .B0 (nx26605), .B1 (
          nx35217)) ;
    aoi32 ix26599 (.Y (nx26598), .A0 (nx5336), .A1 (nx34683), .A2 (nx26603), .B0 (
          mdr_data_out[30]), .B1 (nx34677)) ;
    nand02 ix5337 (.Y (nx5336), .A0 (nx26601), .A1 (mdr_data_out[30])) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_31), .QB (nx26605), .D (nx16903)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix26609 (.Y (nx26608), .A0 (mdr_data_out[31]), .A1 (nx34677), .B0 (
          nx34683), .B1 (nx5356)) ;
    xnor2 ix5357 (.Y (nx5356), .A0 (mdr_data_out[31]), .A1 (nx5340)) ;
    nor02ii ix5341 (.Y (nx5340), .A0 (mdr_data_out[30]), .A1 (nx5316)) ;
    aoi32 ix26613 (.Y (nx26612), .A0 (nx5312), .A1 (nx34683), .A2 (nx26601), .B0 (
          mdr_data_out[29]), .B1 (nx34677)) ;
    aoi32 ix26616 (.Y (nx26615), .A0 (nx5264), .A1 (nx34683), .A2 (nx26566), .B0 (
          mdr_data_out[27]), .B1 (nx34677)) ;
    aoi32 ix26619 (.Y (nx26618), .A0 (nx5216), .A1 (nx34683), .A2 (nx26531), .B0 (
          mdr_data_out[25]), .B1 (nx34677)) ;
    aoi32 ix26622 (.Y (nx26621), .A0 (nx5168), .A1 (nx34683), .A2 (nx26496), .B0 (
          mdr_data_out[23]), .B1 (nx34677)) ;
    aoi32 ix26625 (.Y (nx26624), .A0 (nx5120), .A1 (nx34683), .A2 (nx26461), .B0 (
          mdr_data_out[21]), .B1 (nx34677)) ;
    aoi32 ix26628 (.Y (nx26627), .A0 (nx5072), .A1 (nx5008), .A2 (nx26426), .B0 (
          mdr_data_out[19]), .B1 (nx34679)) ;
    aoi32 ix26631 (.Y (nx26630), .A0 (nx5022), .A1 (nx5008), .A2 (nx26375), .B0 (
          mdr_data_out[17]), .B1 (nx34679)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_0_booth_output_16), .QB (nx26356), .D (nx17043)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_0_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_0_15), .QB (nx26634), .D (nx17053), .CLK (
         clk), .R (rst)) ;
    aoi21 ix5747 (.Y (nx5746), .A0 (label_1_output[0]), .A1 (nx35731), .B0 (
          nx36387)) ;
    dffr reg_sel_dst_0 (.Q (sel_dst_0), .QB (\$dummy [99]), .D (nx14113), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix14114 (.Y (nx14113), .A0 (sel_dst_0), .A1 (nx36201), .S0 (nx878)
             ) ;
    nor03_2x ix879 (.Y (nx878), .A0 (nx12895), .A1 (nx56), .A2 (nx26661)) ;
    oai21 ix26662 (.Y (nx26661), .A0 (nx25944), .A1 (nx35099), .B0 (nx868)) ;
    oai21 ix869 (.Y (nx868), .A0 (nx26664), .A1 (nx26666), .B0 (nx172)) ;
    dff max_calc_reg_ans1_0 (.Q (max_calc_ans1_0), .QB (\$dummy [100]), .D (
        nx17583), .CLK (clk)) ;
    nand04 ix26676 (.Y (nx26675), .A0 (nx25940), .A1 (max_calc_start), .A2 (
           nx26188), .A3 (nx6368)) ;
    aoi21 ix6369 (.Y (nx6368), .A0 (nx35977), .A1 (nx36389), .B0 (
          max_calc_state_3)) ;
    dff max_calc_reg_ans6_0 (.Q (max_calc_ans6_0), .QB (\$dummy [101]), .D (
        nx17593), .CLK (clk)) ;
    dff max_calc_reg_ans5_0 (.Q (max_calc_ans5_0), .QB (\$dummy [102]), .D (
        nx19623), .CLK (clk)) ;
    oai21 ix18154 (.Y (nx18153), .A0 (nx26693), .A1 (nx34747), .B0 (nx26696)) ;
    dff max_calc_reg_comparator_fifth_inp1_0 (.Q (
        max_calc_comparator_fifth_inp1_0), .QB (nx26693), .D (nx18153), .CLK (
        clk)) ;
    nand03 ix26697 (.Y (nx26696), .A0 (label_9_output[0]), .A1 (nx34737), .A2 (
           nx34747)) ;
    dffr labelsregfile_label9_loop1_0_fx_reg_q (.Q (label_9_output[0]), .QB (
         \$dummy [103]), .D (nx18143), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_0 (.Q (label_9_input_0), .D (nx7260), .CLK (nx34511)
          ) ;
    oai21 ix7261 (.Y (nx7260), .A0 (nx26702), .A1 (nx34409), .B0 (nx26706)) ;
    dffr reg_label_9_input_state_machine_0 (.Q (label_9_input_state_machine_0), 
         .QB (nx26702), .D (nx18133), .CLK (clk), .R (rst)) ;
    oai21 ix26707 (.Y (nx26706), .A0 (nx35755), .A1 (label_9_output[0]), .B0 (
          nx7248)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_8_1), .QB (\$dummy [104]), .D (nx18113)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_8_2), .QB (nx27127), .D (nx18103), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_8_3), .QB (\$dummy [105]), .D (nx18093)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_8_4), .QB (nx27125), .D (nx18083), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_8_5), .QB (\$dummy [106]), .D (nx18073)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_8_6), .QB (nx27123), .D (nx18063), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_8_7), .QB (\$dummy [107]), .D (nx18053)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_8_8), .QB (nx27121), .D (nx18043), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_8_9), .QB (\$dummy [108]), .D (nx18033)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_8_10), .QB (nx27119), .D (nx18023), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_8_11), .QB (\$dummy [109]), .D (nx18013)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_8_12), .QB (nx27117), .D (nx18003), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_8_13), .QB (\$dummy [110]), .D (nx17993)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_8_14), .QB (nx27115), .D (nx17983), .CLK (
         clk), .R (rst)) ;
    aoi22 ix26756 (.Y (nx26755), .A0 (mdr_data_out[15]), .A1 (nx34847), .B0 (
          nx7044), .B1 (nx7050)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_reg_output_0), .QB (\$dummy [111]), .D (
         nx17623), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_8_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_8_shift_Reg_count_0), .QB (\$dummy [112]), .D (
            nx17609), .CLK (clk), .S (nx34467)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_reg_output_9), .QB (\$dummy [113]), .D (
         nx17803), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_9), .QB (\$dummy [114]), .D (
         nx17793), .CLK (clk), .R (nx34467)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_8), .QB (\$dummy [115]), .D (
         nx17783), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_8), .QB (\$dummy [116]), .D (
         nx17773), .CLK (clk), .R (nx34467)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_7), .QB (\$dummy [117]), .D (
         nx17763), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_7), .QB (\$dummy [118]), .D (
         nx17753), .CLK (clk), .R (nx34467)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_6), .QB (\$dummy [119]), .D (
         nx17743), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_6), .QB (\$dummy [120]), .D (
         nx17733), .CLK (clk), .R (nx34467)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_5), .QB (\$dummy [121]), .D (
         nx17723), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_5), .QB (\$dummy [122]), .D (
         nx17713), .CLK (clk), .R (nx34467)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_4), .QB (\$dummy [123]), .D (
         nx17703), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_4), .QB (\$dummy [124]), .D (
         nx17693), .CLK (clk), .R (nx34467)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_3), .QB (\$dummy [125]), .D (
         nx17683), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_3), .QB (\$dummy [126]), .D (
         nx17673), .CLK (clk), .R (nx34465)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_2), .QB (\$dummy [127]), .D (
         nx17663), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_2), .QB (\$dummy [128]), .D (
         nx17653), .CLK (clk), .R (nx34465)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_8_shift_Reg_output_1), .QB (\$dummy [129]), .D (
         nx17643), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_8_shift_Reg_count_1), .QB (\$dummy [130]), .D (
         nx17633), .CLK (clk), .R (nx34465)) ;
    nand02 ix17604 (.Y (nx17603), .A0 (nx35807), .A1 (nx34833)) ;
    dffs_ni booth_booth_integrtaion_8_shift_Reg_reg_en (.Q (\$dummy [131]), .QB (
            nx26802), .D (nx17603), .CLK (clk), .S (nx34465)) ;
    nand02 ix7045 (.Y (nx7044), .A0 (nx26823), .A1 (nx26835)) ;
    oai21 ix26824 (.Y (nx26823), .A0 (nx34861), .A1 (nx34855), .B0 (
          mdr_data_out[144])) ;
    oai21 ix17814 (.Y (nx17813), .A0 (nx26828), .A1 (nx35301), .B0 (nx26830)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [132]), .QB (
         nx26828), .D (nx17813), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [133]), .QB (
         nx26832), .D (nx18123), .CLK (clk), .R (rst)) ;
    xnor2 ix26840 (.Y (nx26839), .A0 (nx6514), .A1 (nx13123)) ;
    oai21 ix17954 (.Y (nx17953), .A0 (nx26845), .A1 (nx35301), .B0 (nx26847)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_17), .QB (nx26845), .D (nx17953)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26848 (.Y (nx26847), .A0 (nx35309), .A1 (nx7022), .A2 (nx36031)) ;
    xnor2 ix7023 (.Y (nx7022), .A0 (nx26850), .A1 (nx13125)) ;
    aoi22 ix26851 (.Y (nx26850), .A0 (booth_booth_integrtaion_8_booth_output_17)
          , .A1 (nx6538), .B0 (nx6514), .B1 (nx13123)) ;
    nand02 ix6523 (.Y (nx6522), .A0 (mdr_data_out[145]), .A1 (mdr_data_out[144])
           ) ;
    or02 ix26855 (.Y (nx26854), .A0 (mdr_data_out[144]), .A1 (mdr_data_out[145])
         ) ;
    xnor2 ix26861 (.Y (nx26860), .A0 (nx6566), .A1 (nx13127)) ;
    oai22 ix6567 (.Y (nx6566), .A0 (nx26850), .A1 (nx26863), .B0 (nx26870), .B1 (
          nx35313)) ;
    aoi32 ix26866 (.Y (nx26865), .A0 (nx6548), .A1 (nx34861), .A2 (nx26868), .B0 (
          mdr_data_out[146]), .B1 (nx34855)) ;
    oai21 ix6549 (.Y (nx6548), .A0 (mdr_data_out[144]), .A1 (mdr_data_out[145])
          , .B0 (mdr_data_out[146])) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_18), .QB (nx26870), .D (nx17943)
         , .CLK (clk), .R (rst)) ;
    oai21 ix17934 (.Y (nx17933), .A0 (nx26875), .A1 (nx35301), .B0 (nx26877)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_19), .QB (nx26875), .D (nx17933)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26878 (.Y (nx26877), .A0 (nx35309), .A1 (nx6998), .A2 (nx36031)) ;
    xnor2 ix6999 (.Y (nx6998), .A0 (nx26880), .A1 (nx13129)) ;
    aoi22 ix26881 (.Y (nx26880), .A0 (booth_booth_integrtaion_8_booth_output_19)
          , .A1 (nx6586), .B0 (nx6566), .B1 (nx13127)) ;
    nor02ii ix26884 (.Y (nx26883), .A0 (nx6552), .A1 (mdr_data_out[147])) ;
    nor03_2x ix6553 (.Y (nx6552), .A0 (mdr_data_out[146]), .A1 (
             mdr_data_out[144]), .A2 (mdr_data_out[145])) ;
    nor04 ix6577 (.Y (nx6576), .A0 (mdr_data_out[147]), .A1 (mdr_data_out[146])
          , .A2 (mdr_data_out[144]), .A3 (mdr_data_out[145])) ;
    xnor2 ix26898 (.Y (nx26897), .A0 (nx6614), .A1 (nx13131)) ;
    oai22 ix6615 (.Y (nx6614), .A0 (nx26880), .A1 (nx26900), .B0 (nx26909), .B1 (
          nx35315)) ;
    aoi32 ix26903 (.Y (nx26902), .A0 (nx6596), .A1 (nx34861), .A2 (nx26907), .B0 (
          mdr_data_out[148]), .B1 (nx34855)) ;
    nand02 ix6597 (.Y (nx6596), .A0 (nx26905), .A1 (mdr_data_out[148])) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_20), .QB (nx26909), .D (nx17923)
         , .CLK (clk), .R (rst)) ;
    oai21 ix17914 (.Y (nx17913), .A0 (nx26914), .A1 (nx35301), .B0 (nx26916)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_21), .QB (nx26914), .D (nx17913)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26917 (.Y (nx26916), .A0 (nx35309), .A1 (nx6974), .A2 (nx36031)) ;
    xnor2 ix6975 (.Y (nx6974), .A0 (nx26919), .A1 (nx13133)) ;
    aoi22 ix26920 (.Y (nx26919), .A0 (booth_booth_integrtaion_8_booth_output_21)
          , .A1 (nx6634), .B0 (nx6614), .B1 (nx13131)) ;
    nor02ii ix26923 (.Y (nx26922), .A0 (nx6600), .A1 (mdr_data_out[149])) ;
    nor02ii ix6601 (.Y (nx6600), .A0 (mdr_data_out[148]), .A1 (nx6576)) ;
    nor02ii ix6625 (.Y (nx6624), .A0 (mdr_data_out[149]), .A1 (nx6600)) ;
    xnor2 ix26933 (.Y (nx26932), .A0 (nx6662), .A1 (nx13135)) ;
    oai22 ix6663 (.Y (nx6662), .A0 (nx26919), .A1 (nx26935), .B0 (nx26944), .B1 (
          nx35317)) ;
    aoi32 ix26938 (.Y (nx26937), .A0 (nx6644), .A1 (nx34861), .A2 (nx26942), .B0 (
          mdr_data_out[150]), .B1 (nx34855)) ;
    nand02 ix6645 (.Y (nx6644), .A0 (nx26940), .A1 (mdr_data_out[150])) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_22), .QB (nx26944), .D (nx17903)
         , .CLK (clk), .R (rst)) ;
    oai21 ix17894 (.Y (nx17893), .A0 (nx26949), .A1 (nx35301), .B0 (nx26951)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_23), .QB (nx26949), .D (nx17893)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26952 (.Y (nx26951), .A0 (nx35309), .A1 (nx6950), .A2 (nx35303)) ;
    xnor2 ix6951 (.Y (nx6950), .A0 (nx26954), .A1 (nx13137)) ;
    aoi22 ix26955 (.Y (nx26954), .A0 (booth_booth_integrtaion_8_booth_output_23)
          , .A1 (nx6682), .B0 (nx6662), .B1 (nx13135)) ;
    nor02ii ix26958 (.Y (nx26957), .A0 (nx6648), .A1 (mdr_data_out[151])) ;
    nor02ii ix6649 (.Y (nx6648), .A0 (mdr_data_out[150]), .A1 (nx6624)) ;
    nor02ii ix6673 (.Y (nx6672), .A0 (mdr_data_out[151]), .A1 (nx6648)) ;
    xnor2 ix26968 (.Y (nx26967), .A0 (nx6710), .A1 (nx13138)) ;
    oai22 ix6711 (.Y (nx6710), .A0 (nx26954), .A1 (nx26970), .B0 (nx26979), .B1 (
          nx35319)) ;
    aoi32 ix26973 (.Y (nx26972), .A0 (nx6692), .A1 (nx34861), .A2 (nx26977), .B0 (
          mdr_data_out[152]), .B1 (nx34855)) ;
    nand02 ix6693 (.Y (nx6692), .A0 (nx26975), .A1 (mdr_data_out[152])) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_24), .QB (nx26979), .D (nx17883)
         , .CLK (clk), .R (rst)) ;
    oai21 ix17874 (.Y (nx17873), .A0 (nx26984), .A1 (nx35303), .B0 (nx26986)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_25), .QB (nx26984), .D (nx17873)
         , .CLK (clk), .R (rst)) ;
    nand03 ix26987 (.Y (nx26986), .A0 (nx35309), .A1 (nx6926), .A2 (nx35303)) ;
    xnor2 ix6927 (.Y (nx6926), .A0 (nx26989), .A1 (nx13139)) ;
    aoi22 ix26990 (.Y (nx26989), .A0 (booth_booth_integrtaion_8_booth_output_25)
          , .A1 (nx6730), .B0 (nx6710), .B1 (nx13138)) ;
    nor02ii ix26993 (.Y (nx26992), .A0 (nx6696), .A1 (mdr_data_out[153])) ;
    nor02ii ix6697 (.Y (nx6696), .A0 (mdr_data_out[152]), .A1 (nx6672)) ;
    nor02ii ix6721 (.Y (nx6720), .A0 (mdr_data_out[153]), .A1 (nx6696)) ;
    xnor2 ix27003 (.Y (nx27002), .A0 (nx6758), .A1 (nx13141)) ;
    oai22 ix6759 (.Y (nx6758), .A0 (nx26989), .A1 (nx27005), .B0 (nx27014), .B1 (
          nx35321)) ;
    aoi32 ix27008 (.Y (nx27007), .A0 (nx6740), .A1 (nx34861), .A2 (nx27012), .B0 (
          mdr_data_out[154]), .B1 (nx34855)) ;
    nand02 ix6741 (.Y (nx6740), .A0 (nx27010), .A1 (mdr_data_out[154])) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_26), .QB (nx27014), .D (nx17863)
         , .CLK (clk), .R (rst)) ;
    oai21 ix17854 (.Y (nx17853), .A0 (nx27019), .A1 (nx35303), .B0 (nx27021)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_27), .QB (nx27019), .D (nx17853)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27022 (.Y (nx27021), .A0 (nx35309), .A1 (nx6902), .A2 (nx35303)) ;
    xnor2 ix6903 (.Y (nx6902), .A0 (nx27024), .A1 (nx13143)) ;
    aoi22 ix27025 (.Y (nx27024), .A0 (booth_booth_integrtaion_8_booth_output_27)
          , .A1 (nx6778), .B0 (nx6758), .B1 (nx13141)) ;
    nor02ii ix27028 (.Y (nx27027), .A0 (nx6744), .A1 (mdr_data_out[155])) ;
    nor02ii ix6745 (.Y (nx6744), .A0 (mdr_data_out[154]), .A1 (nx6720)) ;
    nor02ii ix6769 (.Y (nx6768), .A0 (mdr_data_out[155]), .A1 (nx6744)) ;
    xnor2 ix27038 (.Y (nx27037), .A0 (nx6806), .A1 (nx13145)) ;
    oai22 ix6807 (.Y (nx6806), .A0 (nx27024), .A1 (nx27040), .B0 (nx27049), .B1 (
          nx35323)) ;
    aoi32 ix27043 (.Y (nx27042), .A0 (nx6788), .A1 (nx34861), .A2 (nx27047), .B0 (
          mdr_data_out[156]), .B1 (nx34855)) ;
    nand02 ix6789 (.Y (nx6788), .A0 (nx27045), .A1 (mdr_data_out[156])) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_28), .QB (nx27049), .D (nx17843)
         , .CLK (clk), .R (rst)) ;
    oai21 ix17834 (.Y (nx17833), .A0 (nx27054), .A1 (nx35303), .B0 (nx27056)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_29), .QB (nx27054), .D (nx17833)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27057 (.Y (nx27056), .A0 (nx36039), .A1 (nx6878), .A2 (nx35303)) ;
    xnor2 ix6879 (.Y (nx6878), .A0 (nx27059), .A1 (nx13146)) ;
    aoi22 ix27060 (.Y (nx27059), .A0 (booth_booth_integrtaion_8_booth_output_29)
          , .A1 (nx6826), .B0 (nx6806), .B1 (nx13145)) ;
    nor02ii ix27063 (.Y (nx27062), .A0 (nx6792), .A1 (mdr_data_out[157])) ;
    nor02ii ix6793 (.Y (nx6792), .A0 (mdr_data_out[156]), .A1 (nx6768)) ;
    nor02ii ix6817 (.Y (nx6816), .A0 (mdr_data_out[157]), .A1 (nx6792)) ;
    xnor2 ix27073 (.Y (nx27072), .A0 (nx6854), .A1 (nx6864)) ;
    oai22 ix6855 (.Y (nx6854), .A0 (nx27059), .A1 (nx27075), .B0 (nx27084), .B1 (
          nx35325)) ;
    aoi32 ix27078 (.Y (nx27077), .A0 (nx6836), .A1 (nx34863), .A2 (nx27082), .B0 (
          mdr_data_out[158]), .B1 (nx34857)) ;
    nand02 ix6837 (.Y (nx6836), .A0 (nx27080), .A1 (mdr_data_out[158])) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_31), .QB (nx27084), .D (nx17823)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix27088 (.Y (nx27087), .A0 (mdr_data_out[159]), .A1 (nx34857), .B0 (
          nx34863), .B1 (nx6856)) ;
    xnor2 ix6857 (.Y (nx6856), .A0 (mdr_data_out[159]), .A1 (nx6840)) ;
    nor02ii ix6841 (.Y (nx6840), .A0 (mdr_data_out[158]), .A1 (nx6816)) ;
    aoi32 ix27092 (.Y (nx27091), .A0 (nx6812), .A1 (nx34863), .A2 (nx27080), .B0 (
          mdr_data_out[157]), .B1 (nx34857)) ;
    aoi32 ix27095 (.Y (nx27094), .A0 (nx6764), .A1 (nx34863), .A2 (nx27045), .B0 (
          mdr_data_out[155]), .B1 (nx34857)) ;
    aoi32 ix27098 (.Y (nx27097), .A0 (nx6716), .A1 (nx34863), .A2 (nx27010), .B0 (
          mdr_data_out[153]), .B1 (nx34857)) ;
    aoi32 ix27101 (.Y (nx27100), .A0 (nx6668), .A1 (nx34863), .A2 (nx26975), .B0 (
          mdr_data_out[151]), .B1 (nx34857)) ;
    aoi32 ix27104 (.Y (nx27103), .A0 (nx6620), .A1 (nx34863), .A2 (nx26940), .B0 (
          mdr_data_out[149]), .B1 (nx34857)) ;
    aoi32 ix27107 (.Y (nx27106), .A0 (nx6572), .A1 (nx6508), .A2 (nx26905), .B0 (
          mdr_data_out[147]), .B1 (nx34859)) ;
    aoi32 ix27110 (.Y (nx27109), .A0 (nx6522), .A1 (nx6508), .A2 (nx26854), .B0 (
          mdr_data_out[145]), .B1 (nx34859)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_8_booth_output_16), .QB (nx26835), .D (nx17963)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_8_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_8_15), .QB (nx27113), .D (nx17973), .CLK (
         clk), .R (rst)) ;
    aoi21 ix7249 (.Y (nx7248), .A0 (label_9_output[0]), .A1 (nx35755), .B0 (
          nx36387)) ;
    oai21 ix19554 (.Y (nx19553), .A0 (nx27133), .A1 (nx34747), .B0 (nx27135)) ;
    dff max_calc_reg_comparator_fifth_inp2_0 (.Q (\$dummy [134]), .QB (nx27133)
        , .D (nx19553), .CLK (clk)) ;
    nand03 ix27136 (.Y (nx27135), .A0 (label_10_output[0]), .A1 (nx34737), .A2 (
           nx34747)) ;
    dffr labelsregfile_label10_loop1_0_fx_reg_q (.Q (label_10_output[0]), .QB (
         \$dummy [135]), .D (nx18713), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_0 (.Q (label_10_input_0), .D (nx8138), .CLK (
          nx34511)) ;
    oai21 ix8139 (.Y (nx8138), .A0 (nx27141), .A1 (nx34409), .B0 (nx27145)) ;
    dffr reg_label_10_input_state_machine_0 (.Q (label_10_input_state_machine_0)
         , .QB (nx27141), .D (nx18703), .CLK (clk), .R (rst)) ;
    oai21 ix27146 (.Y (nx27145), .A0 (nx35759), .A1 (label_10_output[0]), .B0 (
          nx8126)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_9_1), .QB (\$dummy [136]), .D (nx18683)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_9_2), .QB (nx27566), .D (nx18673), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_9_3), .QB (\$dummy [137]), .D (nx18663)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_9_4), .QB (nx27564), .D (nx18653), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_9_5), .QB (\$dummy [138]), .D (nx18643)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_9_6), .QB (nx27562), .D (nx18633), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_9_7), .QB (\$dummy [139]), .D (nx18623)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_9_8), .QB (nx27560), .D (nx18613), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_9_9), .QB (\$dummy [140]), .D (nx18603)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_9_10), .QB (nx27558), .D (nx18593), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_9_11), .QB (\$dummy [141]), .D (nx18583)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_9_12), .QB (nx27556), .D (nx18573), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_9_13), .QB (\$dummy [142]), .D (nx18563)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_9_14), .QB (nx27554), .D (nx18553), .CLK (
         clk), .R (rst)) ;
    aoi22 ix27195 (.Y (nx27194), .A0 (mdr_data_out[15]), .A1 (nx34879), .B0 (
          nx7924), .B1 (nx7930)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_reg_output_0), .QB (\$dummy [143]), .D (
         nx18193), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_9_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_9_shift_Reg_count_0), .QB (\$dummy [144]), .D (
            nx18179), .CLK (clk), .S (nx34471)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_reg_output_9), .QB (\$dummy [145]), .D (
         nx18373), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_9), .QB (\$dummy [146]), .D (
         nx18363), .CLK (clk), .R (nx34471)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_8), .QB (\$dummy [147]), .D (
         nx18353), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_8), .QB (\$dummy [148]), .D (
         nx18343), .CLK (clk), .R (nx34471)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_7), .QB (\$dummy [149]), .D (
         nx18333), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_7), .QB (\$dummy [150]), .D (
         nx18323), .CLK (clk), .R (nx34471)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_6), .QB (\$dummy [151]), .D (
         nx18313), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_6), .QB (\$dummy [152]), .D (
         nx18303), .CLK (clk), .R (nx34469)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_5), .QB (\$dummy [153]), .D (
         nx18293), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_5), .QB (\$dummy [154]), .D (
         nx18283), .CLK (clk), .R (nx34469)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_4), .QB (\$dummy [155]), .D (
         nx18273), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_4), .QB (\$dummy [156]), .D (
         nx18263), .CLK (clk), .R (nx34469)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_3), .QB (\$dummy [157]), .D (
         nx18253), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_3), .QB (\$dummy [158]), .D (
         nx18243), .CLK (clk), .R (nx34469)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_2), .QB (\$dummy [159]), .D (
         nx18233), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_2), .QB (\$dummy [160]), .D (
         nx18223), .CLK (clk), .R (nx34469)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_9_shift_Reg_output_1), .QB (\$dummy [161]), .D (
         nx18213), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_9_shift_Reg_count_1), .QB (\$dummy [162]), .D (
         nx18203), .CLK (clk), .R (nx34469)) ;
    nand02 ix18174 (.Y (nx18173), .A0 (nx35811), .A1 (nx34865)) ;
    dffs_ni booth_booth_integrtaion_9_shift_Reg_reg_en (.Q (\$dummy [163]), .QB (
            nx27241), .D (nx18173), .CLK (clk), .S (nx34469)) ;
    nand02 ix7925 (.Y (nx7924), .A0 (nx27262), .A1 (nx27274)) ;
    oai21 ix27263 (.Y (nx27262), .A0 (nx34893), .A1 (nx34887), .B0 (
          mdr_data_out[160])) ;
    oai21 ix18384 (.Y (nx18383), .A0 (nx27267), .A1 (nx35327), .B0 (nx27269)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [164]), .QB (
         nx27267), .D (nx18383), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [165]), .QB (
         nx27271), .D (nx18693), .CLK (clk), .R (rst)) ;
    xnor2 ix27279 (.Y (nx27278), .A0 (nx7394), .A1 (nx13149)) ;
    oai21 ix18524 (.Y (nx18523), .A0 (nx27284), .A1 (nx35327), .B0 (nx27286)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_17), .QB (nx27284), .D (nx18523)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27287 (.Y (nx27286), .A0 (nx35335), .A1 (nx7902), .A2 (nx36047)) ;
    xnor2 ix7903 (.Y (nx7902), .A0 (nx27289), .A1 (nx13151)) ;
    aoi22 ix27290 (.Y (nx27289), .A0 (booth_booth_integrtaion_9_booth_output_17)
          , .A1 (nx7418), .B0 (nx7394), .B1 (nx13149)) ;
    nand02 ix7403 (.Y (nx7402), .A0 (mdr_data_out[161]), .A1 (mdr_data_out[160])
           ) ;
    or02 ix27294 (.Y (nx27293), .A0 (mdr_data_out[160]), .A1 (mdr_data_out[161])
         ) ;
    xnor2 ix27300 (.Y (nx27299), .A0 (nx7446), .A1 (nx13153)) ;
    oai22 ix7447 (.Y (nx7446), .A0 (nx27289), .A1 (nx27302), .B0 (nx27309), .B1 (
          nx35339)) ;
    aoi32 ix27305 (.Y (nx27304), .A0 (nx7428), .A1 (nx34893), .A2 (nx27307), .B0 (
          mdr_data_out[162]), .B1 (nx34887)) ;
    oai21 ix7429 (.Y (nx7428), .A0 (mdr_data_out[160]), .A1 (mdr_data_out[161])
          , .B0 (mdr_data_out[162])) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_18), .QB (nx27309), .D (nx18513)
         , .CLK (clk), .R (rst)) ;
    oai21 ix18504 (.Y (nx18503), .A0 (nx27314), .A1 (nx35327), .B0 (nx27316)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_19), .QB (nx27314), .D (nx18503)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27317 (.Y (nx27316), .A0 (nx35335), .A1 (nx7878), .A2 (nx36047)) ;
    xnor2 ix7879 (.Y (nx7878), .A0 (nx27319), .A1 (nx13155)) ;
    aoi22 ix27320 (.Y (nx27319), .A0 (booth_booth_integrtaion_9_booth_output_19)
          , .A1 (nx7466), .B0 (nx7446), .B1 (nx13153)) ;
    nor02ii ix27323 (.Y (nx27322), .A0 (nx7432), .A1 (mdr_data_out[163])) ;
    nor03_2x ix7433 (.Y (nx7432), .A0 (mdr_data_out[162]), .A1 (
             mdr_data_out[160]), .A2 (mdr_data_out[161])) ;
    nor04 ix7457 (.Y (nx7456), .A0 (mdr_data_out[163]), .A1 (mdr_data_out[162])
          , .A2 (mdr_data_out[160]), .A3 (mdr_data_out[161])) ;
    xnor2 ix27337 (.Y (nx27336), .A0 (nx7494), .A1 (nx13157)) ;
    oai22 ix7495 (.Y (nx7494), .A0 (nx27319), .A1 (nx27339), .B0 (nx27348), .B1 (
          nx35341)) ;
    aoi32 ix27342 (.Y (nx27341), .A0 (nx7476), .A1 (nx34893), .A2 (nx27346), .B0 (
          mdr_data_out[164]), .B1 (nx34887)) ;
    nand02 ix7477 (.Y (nx7476), .A0 (nx27344), .A1 (mdr_data_out[164])) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_20), .QB (nx27348), .D (nx18493)
         , .CLK (clk), .R (rst)) ;
    oai21 ix18484 (.Y (nx18483), .A0 (nx27353), .A1 (nx35327), .B0 (nx27355)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_21), .QB (nx27353), .D (nx18483)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27356 (.Y (nx27355), .A0 (nx35335), .A1 (nx7854), .A2 (nx36047)) ;
    xnor2 ix7855 (.Y (nx7854), .A0 (nx27358), .A1 (nx13159)) ;
    aoi22 ix27359 (.Y (nx27358), .A0 (booth_booth_integrtaion_9_booth_output_21)
          , .A1 (nx7514), .B0 (nx7494), .B1 (nx13157)) ;
    nor02ii ix27362 (.Y (nx27361), .A0 (nx7480), .A1 (mdr_data_out[165])) ;
    nor02ii ix7481 (.Y (nx7480), .A0 (mdr_data_out[164]), .A1 (nx7456)) ;
    nor02ii ix7505 (.Y (nx7504), .A0 (mdr_data_out[165]), .A1 (nx7480)) ;
    xnor2 ix27372 (.Y (nx27371), .A0 (nx7542), .A1 (nx13161)) ;
    oai22 ix7543 (.Y (nx7542), .A0 (nx27358), .A1 (nx27374), .B0 (nx27383), .B1 (
          nx35343)) ;
    aoi32 ix27377 (.Y (nx27376), .A0 (nx7524), .A1 (nx34893), .A2 (nx27381), .B0 (
          mdr_data_out[166]), .B1 (nx34887)) ;
    nand02 ix7525 (.Y (nx7524), .A0 (nx27379), .A1 (mdr_data_out[166])) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_22), .QB (nx27383), .D (nx18473)
         , .CLK (clk), .R (rst)) ;
    oai21 ix18464 (.Y (nx18463), .A0 (nx27388), .A1 (nx35327), .B0 (nx27390)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_23), .QB (nx27388), .D (nx18463)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27391 (.Y (nx27390), .A0 (nx35335), .A1 (nx7830), .A2 (nx35329)) ;
    xnor2 ix7831 (.Y (nx7830), .A0 (nx27393), .A1 (nx13162)) ;
    aoi22 ix27394 (.Y (nx27393), .A0 (booth_booth_integrtaion_9_booth_output_23)
          , .A1 (nx7562), .B0 (nx7542), .B1 (nx13161)) ;
    nor02ii ix27397 (.Y (nx27396), .A0 (nx7528), .A1 (mdr_data_out[167])) ;
    nor02ii ix7529 (.Y (nx7528), .A0 (mdr_data_out[166]), .A1 (nx7504)) ;
    nor02ii ix7553 (.Y (nx7552), .A0 (mdr_data_out[167]), .A1 (nx7528)) ;
    xnor2 ix27407 (.Y (nx27406), .A0 (nx7590), .A1 (nx13163)) ;
    oai22 ix7591 (.Y (nx7590), .A0 (nx27393), .A1 (nx27409), .B0 (nx27418), .B1 (
          nx35345)) ;
    aoi32 ix27412 (.Y (nx27411), .A0 (nx7572), .A1 (nx34893), .A2 (nx27416), .B0 (
          mdr_data_out[168]), .B1 (nx34887)) ;
    nand02 ix7573 (.Y (nx7572), .A0 (nx27414), .A1 (mdr_data_out[168])) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_24), .QB (nx27418), .D (nx18453)
         , .CLK (clk), .R (rst)) ;
    oai21 ix18444 (.Y (nx18443), .A0 (nx27423), .A1 (nx35329), .B0 (nx27425)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_25), .QB (nx27423), .D (nx18443)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27426 (.Y (nx27425), .A0 (nx35335), .A1 (nx7806), .A2 (nx35329)) ;
    xnor2 ix7807 (.Y (nx7806), .A0 (nx27428), .A1 (nx13165)) ;
    aoi22 ix27429 (.Y (nx27428), .A0 (booth_booth_integrtaion_9_booth_output_25)
          , .A1 (nx7610), .B0 (nx7590), .B1 (nx13163)) ;
    nor02ii ix27432 (.Y (nx27431), .A0 (nx7576), .A1 (mdr_data_out[169])) ;
    nor02ii ix7577 (.Y (nx7576), .A0 (mdr_data_out[168]), .A1 (nx7552)) ;
    nor02ii ix7601 (.Y (nx7600), .A0 (mdr_data_out[169]), .A1 (nx7576)) ;
    xnor2 ix27442 (.Y (nx27441), .A0 (nx7638), .A1 (nx13167)) ;
    oai22 ix7639 (.Y (nx7638), .A0 (nx27428), .A1 (nx27444), .B0 (nx27453), .B1 (
          nx35347)) ;
    aoi32 ix27447 (.Y (nx27446), .A0 (nx7620), .A1 (nx34893), .A2 (nx27451), .B0 (
          mdr_data_out[170]), .B1 (nx34887)) ;
    nand02 ix7621 (.Y (nx7620), .A0 (nx27449), .A1 (mdr_data_out[170])) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_26), .QB (nx27453), .D (nx18433)
         , .CLK (clk), .R (rst)) ;
    oai21 ix18424 (.Y (nx18423), .A0 (nx27458), .A1 (nx35329), .B0 (nx27460)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_27), .QB (nx27458), .D (nx18423)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27461 (.Y (nx27460), .A0 (nx35335), .A1 (nx7782), .A2 (nx35329)) ;
    xnor2 ix7783 (.Y (nx7782), .A0 (nx27463), .A1 (nx13169)) ;
    aoi22 ix27464 (.Y (nx27463), .A0 (booth_booth_integrtaion_9_booth_output_27)
          , .A1 (nx7658), .B0 (nx7638), .B1 (nx13167)) ;
    nor02ii ix27467 (.Y (nx27466), .A0 (nx7624), .A1 (mdr_data_out[171])) ;
    nor02ii ix7625 (.Y (nx7624), .A0 (mdr_data_out[170]), .A1 (nx7600)) ;
    nor02ii ix7649 (.Y (nx7648), .A0 (mdr_data_out[171]), .A1 (nx7624)) ;
    xnor2 ix27477 (.Y (nx27476), .A0 (nx7686), .A1 (nx13170)) ;
    oai22 ix7687 (.Y (nx7686), .A0 (nx27463), .A1 (nx27479), .B0 (nx27488), .B1 (
          nx35349)) ;
    aoi32 ix27482 (.Y (nx27481), .A0 (nx7668), .A1 (nx34893), .A2 (nx27486), .B0 (
          mdr_data_out[172]), .B1 (nx34887)) ;
    nand02 ix7669 (.Y (nx7668), .A0 (nx27484), .A1 (mdr_data_out[172])) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_28), .QB (nx27488), .D (nx18413)
         , .CLK (clk), .R (rst)) ;
    oai21 ix18404 (.Y (nx18403), .A0 (nx27493), .A1 (nx35329), .B0 (nx27495)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_29), .QB (nx27493), .D (nx18403)
         , .CLK (clk), .R (rst)) ;
    nand03 ix27496 (.Y (nx27495), .A0 (nx36055), .A1 (nx7758), .A2 (nx35329)) ;
    xnor2 ix7759 (.Y (nx7758), .A0 (nx27498), .A1 (nx13171)) ;
    aoi22 ix27499 (.Y (nx27498), .A0 (booth_booth_integrtaion_9_booth_output_29)
          , .A1 (nx7706), .B0 (nx7686), .B1 (nx13170)) ;
    nor02ii ix27502 (.Y (nx27501), .A0 (nx7672), .A1 (mdr_data_out[173])) ;
    nor02ii ix7673 (.Y (nx7672), .A0 (mdr_data_out[172]), .A1 (nx7648)) ;
    nor02ii ix7697 (.Y (nx7696), .A0 (mdr_data_out[173]), .A1 (nx7672)) ;
    xnor2 ix27512 (.Y (nx27511), .A0 (nx7734), .A1 (nx7744)) ;
    oai22 ix7735 (.Y (nx7734), .A0 (nx27498), .A1 (nx27514), .B0 (nx27523), .B1 (
          nx35351)) ;
    aoi32 ix27517 (.Y (nx27516), .A0 (nx7716), .A1 (nx34895), .A2 (nx27521), .B0 (
          mdr_data_out[174]), .B1 (nx34889)) ;
    nand02 ix7717 (.Y (nx7716), .A0 (nx27519), .A1 (mdr_data_out[174])) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_31), .QB (nx27523), .D (nx18393)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix27527 (.Y (nx27526), .A0 (mdr_data_out[175]), .A1 (nx34889), .B0 (
          nx34895), .B1 (nx7736)) ;
    xnor2 ix7737 (.Y (nx7736), .A0 (mdr_data_out[175]), .A1 (nx7720)) ;
    nor02ii ix7721 (.Y (nx7720), .A0 (mdr_data_out[174]), .A1 (nx7696)) ;
    aoi32 ix27531 (.Y (nx27530), .A0 (nx7692), .A1 (nx34895), .A2 (nx27519), .B0 (
          mdr_data_out[173]), .B1 (nx34889)) ;
    aoi32 ix27534 (.Y (nx27533), .A0 (nx7644), .A1 (nx34895), .A2 (nx27484), .B0 (
          mdr_data_out[171]), .B1 (nx34889)) ;
    aoi32 ix27537 (.Y (nx27536), .A0 (nx7596), .A1 (nx34895), .A2 (nx27449), .B0 (
          mdr_data_out[169]), .B1 (nx34889)) ;
    aoi32 ix27540 (.Y (nx27539), .A0 (nx7548), .A1 (nx34895), .A2 (nx27414), .B0 (
          mdr_data_out[167]), .B1 (nx34889)) ;
    aoi32 ix27543 (.Y (nx27542), .A0 (nx7500), .A1 (nx34895), .A2 (nx27379), .B0 (
          mdr_data_out[165]), .B1 (nx34889)) ;
    aoi32 ix27546 (.Y (nx27545), .A0 (nx7452), .A1 (nx7388), .A2 (nx27344), .B0 (
          mdr_data_out[163]), .B1 (nx34891)) ;
    aoi32 ix27549 (.Y (nx27548), .A0 (nx7402), .A1 (nx7388), .A2 (nx27293), .B0 (
          mdr_data_out[161]), .B1 (nx34891)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_9_booth_output_16), .QB (nx27274), .D (nx18533)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_9_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_9_15), .QB (nx27552), .D (nx18543), .CLK (
         clk), .R (rst)) ;
    aoi21 ix8127 (.Y (nx8126), .A0 (label_10_output[0]), .A1 (nx35759), .B0 (
          nx36387)) ;
    xnor2 ix9491 (.Y (nx9490), .A0 (nx27571), .A1 (nx9488)) ;
    aoi22 ix27572 (.Y (nx27571), .A0 (nx27573), .A1 (
          max_calc_comparator_fifth_inp1_14), .B0 (nx9044), .B1 (nx9398)) ;
    dff max_calc_reg_comparator_fifth_inp2_14 (.Q (\$dummy [166]), .QB (nx27573)
        , .D (nx18993), .CLK (clk)) ;
    oai21 ix18994 (.Y (nx18993), .A0 (nx27573), .A1 (nx34747), .B0 (nx27576)) ;
    dffr labelsregfile_label10_loop1_14_fx_reg_q (.Q (label_10_output[14]), .QB (
         nx27760), .D (nx18983), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_14 (.Q (label_10_input_14), .D (nx8574), .CLK (
          nx34515)) ;
    dffr reg_label_10_input_state_machine_14 (.Q (
         label_10_input_state_machine_14), .QB (\$dummy [167]), .D (nx18163), .CLK (
         clk), .R (rst)) ;
    xor2 ix8571 (.Y (nx8570), .A0 (nx27586), .A1 (nx27758)) ;
    aoi22 ix27587 (.Y (nx27586), .A0 (label_10_output[13]), .A1 (
          booth_booth_integration_output_9_13), .B0 (nx8534), .B1 (nx13199)) ;
    dffr labelsregfile_label10_loop1_13_fx_reg_q (.Q (label_10_output[13]), .QB (
         \$dummy [168]), .D (nx18973), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_13 (.Q (label_10_input_13), .D (nx8548), .CLK (
          nx34515)) ;
    dffr reg_label_10_input_state_machine_13 (.Q (
         label_10_input_state_machine_13), .QB (\$dummy [169]), .D (nx18963), .CLK (
         clk), .R (rst)) ;
    xnor2 ix8545 (.Y (nx8544), .A0 (nx8534), .A1 (nx27754)) ;
    oai22 ix8535 (.Y (nx8534), .A0 (nx27597), .A1 (nx27743), .B0 (nx27753), .B1 (
          nx27556)) ;
    aoi22 ix27598 (.Y (nx27597), .A0 (label_10_output[11]), .A1 (
          booth_booth_integration_output_9_11), .B0 (nx8470), .B1 (nx13195)) ;
    dffr labelsregfile_label10_loop1_11_fx_reg_q (.Q (label_10_output[11]), .QB (
         \$dummy [170]), .D (nx18933), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_11 (.Q (label_10_input_11), .D (nx8484), .CLK (
          nx34513)) ;
    dffr reg_label_10_input_state_machine_11 (.Q (
         label_10_input_state_machine_11), .QB (\$dummy [171]), .D (nx18923), .CLK (
         clk), .R (rst)) ;
    xnor2 ix8481 (.Y (nx8480), .A0 (nx8470), .A1 (nx27739)) ;
    oai22 ix8471 (.Y (nx8470), .A0 (nx27608), .A1 (nx27728), .B0 (nx27738), .B1 (
          nx27558)) ;
    aoi22 ix27609 (.Y (nx27608), .A0 (label_10_output[9]), .A1 (
          booth_booth_integration_output_9_9), .B0 (nx8406), .B1 (nx13191)) ;
    dffr labelsregfile_label10_loop1_9_fx_reg_q (.Q (label_10_output[9]), .QB (
         \$dummy [172]), .D (nx18893), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_9 (.Q (label_10_input_9), .D (nx8420), .CLK (
          nx34513)) ;
    dffr reg_label_10_input_state_machine_9 (.Q (label_10_input_state_machine_9)
         , .QB (\$dummy [173]), .D (nx18883), .CLK (clk), .R (rst)) ;
    xnor2 ix8417 (.Y (nx8416), .A0 (nx8406), .A1 (nx27724)) ;
    oai22 ix8407 (.Y (nx8406), .A0 (nx27619), .A1 (nx27713), .B0 (nx27723), .B1 (
          nx27560)) ;
    aoi22 ix27620 (.Y (nx27619), .A0 (label_10_output[7]), .A1 (
          booth_booth_integration_output_9_7), .B0 (nx8342), .B1 (nx13187)) ;
    dffr labelsregfile_label10_loop1_7_fx_reg_q (.Q (label_10_output[7]), .QB (
         \$dummy [174]), .D (nx18853), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_7 (.Q (label_10_input_7), .D (nx8356), .CLK (
          nx34513)) ;
    dffr reg_label_10_input_state_machine_7 (.Q (label_10_input_state_machine_7)
         , .QB (\$dummy [175]), .D (nx18843), .CLK (clk), .R (rst)) ;
    xnor2 ix8353 (.Y (nx8352), .A0 (nx8342), .A1 (nx27709)) ;
    oai22 ix8343 (.Y (nx8342), .A0 (nx27630), .A1 (nx27698), .B0 (nx27708), .B1 (
          nx27562)) ;
    aoi22 ix27631 (.Y (nx27630), .A0 (label_10_output[5]), .A1 (
          booth_booth_integration_output_9_5), .B0 (nx8278), .B1 (nx13183)) ;
    dffr labelsregfile_label10_loop1_5_fx_reg_q (.Q (label_10_output[5]), .QB (
         \$dummy [176]), .D (nx18813), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_5 (.Q (label_10_input_5), .D (nx8292), .CLK (
          nx34513)) ;
    dffr reg_label_10_input_state_machine_5 (.Q (label_10_input_state_machine_5)
         , .QB (\$dummy [177]), .D (nx18803), .CLK (clk), .R (rst)) ;
    xnor2 ix8289 (.Y (nx8288), .A0 (nx8278), .A1 (nx27694)) ;
    oai22 ix8279 (.Y (nx8278), .A0 (nx27641), .A1 (nx27683), .B0 (nx27693), .B1 (
          nx27564)) ;
    aoi22 ix27642 (.Y (nx27641), .A0 (label_10_output[3]), .A1 (
          booth_booth_integration_output_9_3), .B0 (nx8214), .B1 (nx13179)) ;
    dffr labelsregfile_label10_loop1_3_fx_reg_q (.Q (label_10_output[3]), .QB (
         \$dummy [178]), .D (nx18773), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_3 (.Q (label_10_input_3), .D (nx8228), .CLK (
          nx34511)) ;
    dffr reg_label_10_input_state_machine_3 (.Q (label_10_input_state_machine_3)
         , .QB (\$dummy [179]), .D (nx18763), .CLK (clk), .R (rst)) ;
    xnor2 ix8225 (.Y (nx8224), .A0 (nx8214), .A1 (nx27679)) ;
    oai22 ix8215 (.Y (nx8214), .A0 (nx27652), .A1 (nx27668), .B0 (nx27678), .B1 (
          nx27566)) ;
    aoi32 ix27653 (.Y (nx27652), .A0 (label_10_output[0]), .A1 (nx35759), .A2 (
          nx13175), .B0 (label_10_output[1]), .B1 (
          booth_booth_integration_output_9_1)) ;
    dffr labelsregfile_label10_loop1_1_fx_reg_q (.Q (label_10_output[1]), .QB (
         \$dummy [180]), .D (nx18733), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_1 (.Q (label_10_input_1), .D (nx8164), .CLK (
          nx34511)) ;
    dffr reg_label_10_input_state_machine_1 (.Q (label_10_input_state_machine_1)
         , .QB (\$dummy [181]), .D (nx18723), .CLK (clk), .R (rst)) ;
    xor2 ix8161 (.Y (nx8160), .A0 (nx27663), .A1 (nx27665)) ;
    nand02 ix27664 (.Y (nx27663), .A0 (label_10_output[0]), .A1 (nx35759)) ;
    xnor2 ix27666 (.Y (nx27665), .A0 (booth_booth_integration_output_9_1), .A1 (
          label_10_output[1])) ;
    dffr labelsregfile_label10_loop1_2_fx_reg_q (.Q (label_10_output[2]), .QB (
         nx27678), .D (nx18753), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_2 (.Q (label_10_input_2), .D (nx8196), .CLK (
          nx34511)) ;
    dffr reg_label_10_input_state_machine_2 (.Q (label_10_input_state_machine_2)
         , .QB (\$dummy [182]), .D (nx18743), .CLK (clk), .R (rst)) ;
    xor2 ix8193 (.Y (nx8192), .A0 (nx27652), .A1 (nx27668)) ;
    xnor2 ix27680 (.Y (nx27679), .A0 (booth_booth_integration_output_9_3), .A1 (
          label_10_output[3])) ;
    dffr labelsregfile_label10_loop1_4_fx_reg_q (.Q (label_10_output[4]), .QB (
         nx27693), .D (nx18793), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_4 (.Q (label_10_input_4), .D (nx8260), .CLK (
          nx34511)) ;
    dffr reg_label_10_input_state_machine_4 (.Q (label_10_input_state_machine_4)
         , .QB (\$dummy [183]), .D (nx18783), .CLK (clk), .R (rst)) ;
    xor2 ix8257 (.Y (nx8256), .A0 (nx27641), .A1 (nx27683)) ;
    xnor2 ix27695 (.Y (nx27694), .A0 (booth_booth_integration_output_9_5), .A1 (
          label_10_output[5])) ;
    dffr labelsregfile_label10_loop1_6_fx_reg_q (.Q (label_10_output[6]), .QB (
         nx27708), .D (nx18833), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_6 (.Q (label_10_input_6), .D (nx8324), .CLK (
          nx34513)) ;
    dffr reg_label_10_input_state_machine_6 (.Q (label_10_input_state_machine_6)
         , .QB (\$dummy [184]), .D (nx18823), .CLK (clk), .R (rst)) ;
    xor2 ix8321 (.Y (nx8320), .A0 (nx27630), .A1 (nx27698)) ;
    xnor2 ix27710 (.Y (nx27709), .A0 (booth_booth_integration_output_9_7), .A1 (
          label_10_output[7])) ;
    dffr labelsregfile_label10_loop1_8_fx_reg_q (.Q (label_10_output[8]), .QB (
         nx27723), .D (nx18873), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_8 (.Q (label_10_input_8), .D (nx8388), .CLK (
          nx34513)) ;
    dffr reg_label_10_input_state_machine_8 (.Q (label_10_input_state_machine_8)
         , .QB (\$dummy [185]), .D (nx18863), .CLK (clk), .R (rst)) ;
    xor2 ix8385 (.Y (nx8384), .A0 (nx27619), .A1 (nx27713)) ;
    xnor2 ix27725 (.Y (nx27724), .A0 (booth_booth_integration_output_9_9), .A1 (
          label_10_output[9])) ;
    dffr labelsregfile_label10_loop1_10_fx_reg_q (.Q (label_10_output[10]), .QB (
         nx27738), .D (nx18913), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_10 (.Q (label_10_input_10), .D (nx8452), .CLK (
          nx34513)) ;
    dffr reg_label_10_input_state_machine_10 (.Q (
         label_10_input_state_machine_10), .QB (\$dummy [186]), .D (nx18903), .CLK (
         clk), .R (rst)) ;
    xor2 ix8449 (.Y (nx8448), .A0 (nx27608), .A1 (nx27728)) ;
    xnor2 ix27740 (.Y (nx27739), .A0 (booth_booth_integration_output_9_11), .A1 (
          label_10_output[11])) ;
    dffr labelsregfile_label10_loop1_12_fx_reg_q (.Q (label_10_output[12]), .QB (
         nx27753), .D (nx18953), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_12 (.Q (label_10_input_12), .D (nx8516), .CLK (
          nx34515)) ;
    dffr reg_label_10_input_state_machine_12 (.Q (
         label_10_input_state_machine_12), .QB (\$dummy [187]), .D (nx18943), .CLK (
         clk), .R (rst)) ;
    xor2 ix8513 (.Y (nx8512), .A0 (nx27597), .A1 (nx27743)) ;
    xnor2 ix27755 (.Y (nx27754), .A0 (booth_booth_integration_output_9_13), .A1 (
          label_10_output[13])) ;
    oai21 ix19284 (.Y (nx19283), .A0 (nx27763), .A1 (nx34747), .B0 (nx27765)) ;
    dff max_calc_reg_comparator_fifth_inp1_14 (.Q (
        max_calc_comparator_fifth_inp1_14), .QB (nx27763), .D (nx19283), .CLK (
        clk)) ;
    dffr labelsregfile_label9_loop1_14_fx_reg_q (.Q (label_9_output[14]), .QB (
         nx27949), .D (nx19273), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_14 (.Q (label_9_input_14), .D (nx9024), .CLK (
          nx34519)) ;
    dffr reg_label_9_input_state_machine_14 (.Q (label_9_input_state_machine_14)
         , .QB (\$dummy [188]), .D (nx19003), .CLK (clk), .R (rst)) ;
    xor2 ix9021 (.Y (nx9020), .A0 (nx27775), .A1 (nx27947)) ;
    aoi22 ix27776 (.Y (nx27775), .A0 (label_9_output[13]), .A1 (
          booth_booth_integration_output_8_13), .B0 (nx8984), .B1 (nx13215)) ;
    dffr labelsregfile_label9_loop1_13_fx_reg_q (.Q (label_9_output[13]), .QB (
         \$dummy [189]), .D (nx19263), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_13 (.Q (label_9_input_13), .D (nx8998), .CLK (
          nx34519)) ;
    dffr reg_label_9_input_state_machine_13 (.Q (label_9_input_state_machine_13)
         , .QB (\$dummy [190]), .D (nx19253), .CLK (clk), .R (rst)) ;
    xnor2 ix8995 (.Y (nx8994), .A0 (nx8984), .A1 (nx27943)) ;
    oai22 ix8985 (.Y (nx8984), .A0 (nx27786), .A1 (nx27932), .B0 (nx27942), .B1 (
          nx27117)) ;
    aoi22 ix27787 (.Y (nx27786), .A0 (label_9_output[11]), .A1 (
          booth_booth_integration_output_8_11), .B0 (nx8920), .B1 (nx13213)) ;
    dffr labelsregfile_label9_loop1_11_fx_reg_q (.Q (label_9_output[11]), .QB (
         \$dummy [191]), .D (nx19223), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_11 (.Q (label_9_input_11), .D (nx8934), .CLK (
          nx34517)) ;
    dffr reg_label_9_input_state_machine_11 (.Q (label_9_input_state_machine_11)
         , .QB (\$dummy [192]), .D (nx19213), .CLK (clk), .R (rst)) ;
    xnor2 ix8931 (.Y (nx8930), .A0 (nx8920), .A1 (nx27928)) ;
    oai22 ix8921 (.Y (nx8920), .A0 (nx27797), .A1 (nx27917), .B0 (nx27927), .B1 (
          nx27119)) ;
    aoi22 ix27798 (.Y (nx27797), .A0 (label_9_output[9]), .A1 (
          booth_booth_integration_output_8_9), .B0 (nx8856), .B1 (nx13211)) ;
    dffr labelsregfile_label9_loop1_9_fx_reg_q (.Q (label_9_output[9]), .QB (
         \$dummy [193]), .D (nx19183), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_9 (.Q (label_9_input_9), .D (nx8870), .CLK (nx34517)
          ) ;
    dffr reg_label_9_input_state_machine_9 (.Q (label_9_input_state_machine_9), 
         .QB (\$dummy [194]), .D (nx19173), .CLK (clk), .R (rst)) ;
    xnor2 ix8867 (.Y (nx8866), .A0 (nx8856), .A1 (nx27913)) ;
    oai22 ix8857 (.Y (nx8856), .A0 (nx27808), .A1 (nx27902), .B0 (nx27912), .B1 (
          nx27121)) ;
    aoi22 ix27809 (.Y (nx27808), .A0 (label_9_output[7]), .A1 (
          booth_booth_integration_output_8_7), .B0 (nx8792), .B1 (nx13207)) ;
    dffr labelsregfile_label9_loop1_7_fx_reg_q (.Q (label_9_output[7]), .QB (
         \$dummy [195]), .D (nx19143), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_7 (.Q (label_9_input_7), .D (nx8806), .CLK (nx34517)
          ) ;
    dffr reg_label_9_input_state_machine_7 (.Q (label_9_input_state_machine_7), 
         .QB (\$dummy [196]), .D (nx19133), .CLK (clk), .R (rst)) ;
    xnor2 ix8803 (.Y (nx8802), .A0 (nx8792), .A1 (nx27898)) ;
    oai22 ix8793 (.Y (nx8792), .A0 (nx27819), .A1 (nx27887), .B0 (nx27897), .B1 (
          nx27123)) ;
    aoi22 ix27820 (.Y (nx27819), .A0 (label_9_output[5]), .A1 (
          booth_booth_integration_output_8_5), .B0 (nx8728), .B1 (nx13204)) ;
    dffr labelsregfile_label9_loop1_5_fx_reg_q (.Q (label_9_output[5]), .QB (
         \$dummy [197]), .D (nx19103), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_5 (.Q (label_9_input_5), .D (nx8742), .CLK (nx34517)
          ) ;
    dffr reg_label_9_input_state_machine_5 (.Q (label_9_input_state_machine_5), 
         .QB (\$dummy [198]), .D (nx19093), .CLK (clk), .R (rst)) ;
    xnor2 ix8739 (.Y (nx8738), .A0 (nx8728), .A1 (nx27883)) ;
    oai22 ix8729 (.Y (nx8728), .A0 (nx27830), .A1 (nx27872), .B0 (nx27882), .B1 (
          nx27125)) ;
    aoi22 ix27831 (.Y (nx27830), .A0 (label_9_output[3]), .A1 (
          booth_booth_integration_output_8_3), .B0 (nx8664), .B1 (nx13202)) ;
    dffr labelsregfile_label9_loop1_3_fx_reg_q (.Q (label_9_output[3]), .QB (
         \$dummy [199]), .D (nx19063), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_3 (.Q (label_9_input_3), .D (nx8678), .CLK (nx34515)
          ) ;
    dffr reg_label_9_input_state_machine_3 (.Q (label_9_input_state_machine_3), 
         .QB (\$dummy [200]), .D (nx19053), .CLK (clk), .R (rst)) ;
    xnor2 ix8675 (.Y (nx8674), .A0 (nx8664), .A1 (nx27868)) ;
    oai22 ix8665 (.Y (nx8664), .A0 (nx27841), .A1 (nx27857), .B0 (nx27867), .B1 (
          nx27127)) ;
    aoi32 ix27842 (.Y (nx27841), .A0 (label_9_output[0]), .A1 (nx35755), .A2 (
          nx13200), .B0 (label_9_output[1]), .B1 (
          booth_booth_integration_output_8_1)) ;
    dffr labelsregfile_label9_loop1_1_fx_reg_q (.Q (label_9_output[1]), .QB (
         \$dummy [201]), .D (nx19023), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_1 (.Q (label_9_input_1), .D (nx8614), .CLK (nx34515)
          ) ;
    dffr reg_label_9_input_state_machine_1 (.Q (label_9_input_state_machine_1), 
         .QB (\$dummy [202]), .D (nx19013), .CLK (clk), .R (rst)) ;
    xor2 ix8611 (.Y (nx8610), .A0 (nx27852), .A1 (nx27854)) ;
    nand02 ix27853 (.Y (nx27852), .A0 (label_9_output[0]), .A1 (nx35755)) ;
    xnor2 ix27855 (.Y (nx27854), .A0 (booth_booth_integration_output_8_1), .A1 (
          label_9_output[1])) ;
    dffr labelsregfile_label9_loop1_2_fx_reg_q (.Q (label_9_output[2]), .QB (
         nx27867), .D (nx19043), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_2 (.Q (label_9_input_2), .D (nx8646), .CLK (nx34515)
          ) ;
    dffr reg_label_9_input_state_machine_2 (.Q (label_9_input_state_machine_2), 
         .QB (\$dummy [203]), .D (nx19033), .CLK (clk), .R (rst)) ;
    xor2 ix8643 (.Y (nx8642), .A0 (nx27841), .A1 (nx27857)) ;
    xnor2 ix27869 (.Y (nx27868), .A0 (booth_booth_integration_output_8_3), .A1 (
          label_9_output[3])) ;
    dffr labelsregfile_label9_loop1_4_fx_reg_q (.Q (label_9_output[4]), .QB (
         nx27882), .D (nx19083), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_4 (.Q (label_9_input_4), .D (nx8710), .CLK (nx34515)
          ) ;
    dffr reg_label_9_input_state_machine_4 (.Q (label_9_input_state_machine_4), 
         .QB (\$dummy [204]), .D (nx19073), .CLK (clk), .R (rst)) ;
    xor2 ix8707 (.Y (nx8706), .A0 (nx27830), .A1 (nx27872)) ;
    xnor2 ix27884 (.Y (nx27883), .A0 (booth_booth_integration_output_8_5), .A1 (
          label_9_output[5])) ;
    dffr labelsregfile_label9_loop1_6_fx_reg_q (.Q (label_9_output[6]), .QB (
         nx27897), .D (nx19123), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_6 (.Q (label_9_input_6), .D (nx8774), .CLK (nx34517)
          ) ;
    dffr reg_label_9_input_state_machine_6 (.Q (label_9_input_state_machine_6), 
         .QB (\$dummy [205]), .D (nx19113), .CLK (clk), .R (rst)) ;
    xor2 ix8771 (.Y (nx8770), .A0 (nx27819), .A1 (nx27887)) ;
    xnor2 ix27899 (.Y (nx27898), .A0 (booth_booth_integration_output_8_7), .A1 (
          label_9_output[7])) ;
    dffr labelsregfile_label9_loop1_8_fx_reg_q (.Q (label_9_output[8]), .QB (
         nx27912), .D (nx19163), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_8 (.Q (label_9_input_8), .D (nx8838), .CLK (nx34517)
          ) ;
    dffr reg_label_9_input_state_machine_8 (.Q (label_9_input_state_machine_8), 
         .QB (\$dummy [206]), .D (nx19153), .CLK (clk), .R (rst)) ;
    xor2 ix8835 (.Y (nx8834), .A0 (nx27808), .A1 (nx27902)) ;
    xnor2 ix27914 (.Y (nx27913), .A0 (booth_booth_integration_output_8_9), .A1 (
          label_9_output[9])) ;
    dffr labelsregfile_label9_loop1_10_fx_reg_q (.Q (label_9_output[10]), .QB (
         nx27927), .D (nx19203), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_10 (.Q (label_9_input_10), .D (nx8902), .CLK (
          nx34517)) ;
    dffr reg_label_9_input_state_machine_10 (.Q (label_9_input_state_machine_10)
         , .QB (\$dummy [207]), .D (nx19193), .CLK (clk), .R (rst)) ;
    xor2 ix8899 (.Y (nx8898), .A0 (nx27797), .A1 (nx27917)) ;
    xnor2 ix27929 (.Y (nx27928), .A0 (booth_booth_integration_output_8_11), .A1 (
          label_9_output[11])) ;
    dffr labelsregfile_label9_loop1_12_fx_reg_q (.Q (label_9_output[12]), .QB (
         nx27942), .D (nx19243), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_12 (.Q (label_9_input_12), .D (nx8966), .CLK (
          nx34519)) ;
    dffr reg_label_9_input_state_machine_12 (.Q (label_9_input_state_machine_12)
         , .QB (\$dummy [208]), .D (nx19233), .CLK (clk), .R (rst)) ;
    xor2 ix8963 (.Y (nx8962), .A0 (nx27786), .A1 (nx27932)) ;
    xnor2 ix27944 (.Y (nx27943), .A0 (booth_booth_integration_output_8_13), .A1 (
          label_9_output[13])) ;
    oai22 ix9399 (.Y (nx9398), .A0 (nx27952), .A1 (nx27965), .B0 (
          max_calc_comparator_fifth_inp2_13), .B1 (nx27960)) ;
    oai21 ix19294 (.Y (nx19293), .A0 (nx27956), .A1 (nx34749), .B0 (nx27958)) ;
    dff max_calc_reg_comparator_fifth_inp2_13 (.Q (
        max_calc_comparator_fifth_inp2_13), .QB (nx27956), .D (nx19293), .CLK (
        clk)) ;
    nand03 ix27959 (.Y (nx27958), .A0 (label_10_output[13]), .A1 (nx34737), .A2 (
           nx34749)) ;
    dff max_calc_reg_comparator_fifth_inp1_13 (.Q (
        max_calc_comparator_fifth_inp1_13), .QB (nx27960), .D (nx19303), .CLK (
        clk)) ;
    oai21 ix19304 (.Y (nx19303), .A0 (nx27960), .A1 (nx34749), .B0 (nx27963)) ;
    nand03 ix27964 (.Y (nx27963), .A0 (label_9_output[13]), .A1 (nx34739), .A2 (
           nx34749)) ;
    aoi22 ix27966 (.Y (nx27965), .A0 (nx27967), .A1 (
          max_calc_comparator_fifth_inp1_12), .B0 (nx9080), .B1 (nx9382)) ;
    dff max_calc_reg_comparator_fifth_inp2_12 (.Q (\$dummy [209]), .QB (nx27967)
        , .D (nx19313), .CLK (clk)) ;
    oai21 ix19314 (.Y (nx19313), .A0 (nx27967), .A1 (nx34749), .B0 (nx27970)) ;
    oai21 ix19324 (.Y (nx19323), .A0 (nx27974), .A1 (nx34751), .B0 (nx27976)) ;
    dff max_calc_reg_comparator_fifth_inp1_12 (.Q (
        max_calc_comparator_fifth_inp1_12), .QB (nx27974), .D (nx19323), .CLK (
        clk)) ;
    oai22 ix9383 (.Y (nx9382), .A0 (nx27980), .A1 (nx27993), .B0 (
          max_calc_comparator_fifth_inp2_11), .B1 (nx27988)) ;
    oai21 ix19334 (.Y (nx19333), .A0 (nx27984), .A1 (nx34751), .B0 (nx27986)) ;
    dff max_calc_reg_comparator_fifth_inp2_11 (.Q (
        max_calc_comparator_fifth_inp2_11), .QB (nx27984), .D (nx19333), .CLK (
        clk)) ;
    nand03 ix27987 (.Y (nx27986), .A0 (label_10_output[11]), .A1 (nx34739), .A2 (
           nx34751)) ;
    dff max_calc_reg_comparator_fifth_inp1_11 (.Q (
        max_calc_comparator_fifth_inp1_11), .QB (nx27988), .D (nx19343), .CLK (
        clk)) ;
    oai21 ix19344 (.Y (nx19343), .A0 (nx27988), .A1 (nx34751), .B0 (nx27991)) ;
    nand03 ix27992 (.Y (nx27991), .A0 (label_9_output[11]), .A1 (nx34739), .A2 (
           nx34751)) ;
    aoi22 ix27994 (.Y (nx27993), .A0 (nx27995), .A1 (
          max_calc_comparator_fifth_inp1_10), .B0 (nx9116), .B1 (nx9366)) ;
    dff max_calc_reg_comparator_fifth_inp2_10 (.Q (\$dummy [210]), .QB (nx27995)
        , .D (nx19353), .CLK (clk)) ;
    oai21 ix19354 (.Y (nx19353), .A0 (nx27995), .A1 (nx34751), .B0 (nx27998)) ;
    oai21 ix19364 (.Y (nx19363), .A0 (nx28002), .A1 (nx34753), .B0 (nx28004)) ;
    dff max_calc_reg_comparator_fifth_inp1_10 (.Q (
        max_calc_comparator_fifth_inp1_10), .QB (nx28002), .D (nx19363), .CLK (
        clk)) ;
    oai22 ix9367 (.Y (nx9366), .A0 (nx28008), .A1 (nx28021), .B0 (
          max_calc_comparator_fifth_inp2_9), .B1 (nx28016)) ;
    oai21 ix19374 (.Y (nx19373), .A0 (nx28012), .A1 (nx34753), .B0 (nx28014)) ;
    dff max_calc_reg_comparator_fifth_inp2_9 (.Q (
        max_calc_comparator_fifth_inp2_9), .QB (nx28012), .D (nx19373), .CLK (
        clk)) ;
    nand03 ix28015 (.Y (nx28014), .A0 (label_10_output[9]), .A1 (nx34741), .A2 (
           nx34753)) ;
    dff max_calc_reg_comparator_fifth_inp1_9 (.Q (
        max_calc_comparator_fifth_inp1_9), .QB (nx28016), .D (nx19383), .CLK (
        clk)) ;
    oai21 ix19384 (.Y (nx19383), .A0 (nx28016), .A1 (nx34753), .B0 (nx28019)) ;
    nand03 ix28020 (.Y (nx28019), .A0 (label_9_output[9]), .A1 (nx34741), .A2 (
           nx34753)) ;
    aoi22 ix28022 (.Y (nx28021), .A0 (nx28023), .A1 (
          max_calc_comparator_fifth_inp1_8), .B0 (nx9152), .B1 (nx9350)) ;
    dff max_calc_reg_comparator_fifth_inp2_8 (.Q (\$dummy [211]), .QB (nx28023)
        , .D (nx19393), .CLK (clk)) ;
    oai21 ix19394 (.Y (nx19393), .A0 (nx28023), .A1 (nx34755), .B0 (nx28026)) ;
    oai21 ix19404 (.Y (nx19403), .A0 (nx28030), .A1 (nx34755), .B0 (nx28032)) ;
    dff max_calc_reg_comparator_fifth_inp1_8 (.Q (
        max_calc_comparator_fifth_inp1_8), .QB (nx28030), .D (nx19403), .CLK (
        clk)) ;
    oai22 ix9351 (.Y (nx9350), .A0 (nx28036), .A1 (nx28049), .B0 (
          max_calc_comparator_fifth_inp2_7), .B1 (nx28044)) ;
    oai21 ix19414 (.Y (nx19413), .A0 (nx28040), .A1 (nx34755), .B0 (nx28042)) ;
    dff max_calc_reg_comparator_fifth_inp2_7 (.Q (
        max_calc_comparator_fifth_inp2_7), .QB (nx28040), .D (nx19413), .CLK (
        clk)) ;
    nand03 ix28043 (.Y (nx28042), .A0 (label_10_output[7]), .A1 (nx34741), .A2 (
           nx34755)) ;
    dff max_calc_reg_comparator_fifth_inp1_7 (.Q (
        max_calc_comparator_fifth_inp1_7), .QB (nx28044), .D (nx19423), .CLK (
        clk)) ;
    oai21 ix19424 (.Y (nx19423), .A0 (nx28044), .A1 (nx34755), .B0 (nx28047)) ;
    nand03 ix28048 (.Y (nx28047), .A0 (label_9_output[7]), .A1 (nx34741), .A2 (
           nx34757)) ;
    aoi22 ix28050 (.Y (nx28049), .A0 (nx28051), .A1 (
          max_calc_comparator_fifth_inp1_6), .B0 (nx9188), .B1 (nx9334)) ;
    dff max_calc_reg_comparator_fifth_inp2_6 (.Q (\$dummy [212]), .QB (nx28051)
        , .D (nx19433), .CLK (clk)) ;
    oai21 ix19434 (.Y (nx19433), .A0 (nx28051), .A1 (nx34757), .B0 (nx28054)) ;
    oai21 ix19444 (.Y (nx19443), .A0 (nx28058), .A1 (nx34757), .B0 (nx28060)) ;
    dff max_calc_reg_comparator_fifth_inp1_6 (.Q (
        max_calc_comparator_fifth_inp1_6), .QB (nx28058), .D (nx19443), .CLK (
        clk)) ;
    oai22 ix9335 (.Y (nx9334), .A0 (nx28064), .A1 (nx28077), .B0 (
          max_calc_comparator_fifth_inp2_5), .B1 (nx28072)) ;
    oai21 ix19454 (.Y (nx19453), .A0 (nx28068), .A1 (nx34757), .B0 (nx28070)) ;
    dff max_calc_reg_comparator_fifth_inp2_5 (.Q (
        max_calc_comparator_fifth_inp2_5), .QB (nx28068), .D (nx19453), .CLK (
        clk)) ;
    nand03 ix28071 (.Y (nx28070), .A0 (label_10_output[5]), .A1 (nx34743), .A2 (
           nx34757)) ;
    dff max_calc_reg_comparator_fifth_inp1_5 (.Q (
        max_calc_comparator_fifth_inp1_5), .QB (nx28072), .D (nx19463), .CLK (
        clk)) ;
    oai21 ix19464 (.Y (nx19463), .A0 (nx28072), .A1 (nx34759), .B0 (nx28075)) ;
    nand03 ix28076 (.Y (nx28075), .A0 (label_9_output[5]), .A1 (nx34743), .A2 (
           nx34759)) ;
    aoi22 ix28078 (.Y (nx28077), .A0 (nx28079), .A1 (
          max_calc_comparator_fifth_inp1_4), .B0 (nx9224), .B1 (nx9318)) ;
    dff max_calc_reg_comparator_fifth_inp2_4 (.Q (\$dummy [213]), .QB (nx28079)
        , .D (nx19473), .CLK (clk)) ;
    oai21 ix19474 (.Y (nx19473), .A0 (nx28079), .A1 (nx34759), .B0 (nx28082)) ;
    oai21 ix19484 (.Y (nx19483), .A0 (nx28086), .A1 (nx34759), .B0 (nx28088)) ;
    dff max_calc_reg_comparator_fifth_inp1_4 (.Q (
        max_calc_comparator_fifth_inp1_4), .QB (nx28086), .D (nx19483), .CLK (
        clk)) ;
    oai22 ix9319 (.Y (nx9318), .A0 (nx28092), .A1 (nx28105), .B0 (
          max_calc_comparator_fifth_inp2_3), .B1 (nx28100)) ;
    oai21 ix19494 (.Y (nx19493), .A0 (nx28096), .A1 (nx34759), .B0 (nx28098)) ;
    dff max_calc_reg_comparator_fifth_inp2_3 (.Q (
        max_calc_comparator_fifth_inp2_3), .QB (nx28096), .D (nx19493), .CLK (
        clk)) ;
    nand03 ix28099 (.Y (nx28098), .A0 (label_10_output[3]), .A1 (nx34743), .A2 (
           nx34761)) ;
    dff max_calc_reg_comparator_fifth_inp1_3 (.Q (
        max_calc_comparator_fifth_inp1_3), .QB (nx28100), .D (nx19503), .CLK (
        clk)) ;
    oai21 ix19504 (.Y (nx19503), .A0 (nx28100), .A1 (nx34761), .B0 (nx28103)) ;
    nand03 ix28104 (.Y (nx28103), .A0 (label_9_output[3]), .A1 (nx34743), .A2 (
           nx34761)) ;
    aoi22 ix28106 (.Y (nx28105), .A0 (nx28107), .A1 (
          max_calc_comparator_fifth_inp1_2), .B0 (nx9260), .B1 (nx9302)) ;
    dff max_calc_reg_comparator_fifth_inp2_2 (.Q (\$dummy [214]), .QB (nx28107)
        , .D (nx19513), .CLK (clk)) ;
    oai21 ix19514 (.Y (nx19513), .A0 (nx28107), .A1 (nx34761), .B0 (nx28110)) ;
    oai21 ix19524 (.Y (nx19523), .A0 (nx28114), .A1 (nx34761), .B0 (nx28116)) ;
    dff max_calc_reg_comparator_fifth_inp1_2 (.Q (
        max_calc_comparator_fifth_inp1_2), .QB (nx28114), .D (nx19523), .CLK (
        clk)) ;
    oai21 ix9303 (.Y (nx9302), .A0 (max_calc_comparator_fifth_inp2_1), .A1 (
          nx28126), .B0 (nx28131)) ;
    oai21 ix19534 (.Y (nx19533), .A0 (nx28122), .A1 (nx34763), .B0 (nx28124)) ;
    dff max_calc_reg_comparator_fifth_inp2_1 (.Q (
        max_calc_comparator_fifth_inp2_1), .QB (nx28122), .D (nx19533), .CLK (
        clk)) ;
    nand03 ix28125 (.Y (nx28124), .A0 (label_10_output[1]), .A1 (nx34745), .A2 (
           nx34763)) ;
    dff max_calc_reg_comparator_fifth_inp1_1 (.Q (\$dummy [215]), .QB (nx28126)
        , .D (nx19543), .CLK (clk)) ;
    oai21 ix19544 (.Y (nx19543), .A0 (nx28126), .A1 (nx34763), .B0 (nx28129)) ;
    nand03 ix28130 (.Y (nx28129), .A0 (label_9_output[1]), .A1 (nx34745), .A2 (
           nx34763)) ;
    oai21 ix28132 (.Y (nx28131), .A0 (nx27133), .A1 (
          max_calc_comparator_fifth_inp1_0), .B0 (nx9278)) ;
    oai21 ix19584 (.Y (nx19583), .A0 (nx28137), .A1 (nx34763), .B0 (nx28139)) ;
    dff max_calc_reg_comparator_fifth_inp2_15 (.Q (\$dummy [216]), .QB (nx28137)
        , .D (nx19583), .CLK (clk)) ;
    nand03 ix28140 (.Y (nx28139), .A0 (label_10_output[15]), .A1 (nx34745), .A2 (
           nx34763)) ;
    dffr labelsregfile_label10_loop1_15_fx_reg_q (.Q (label_10_output[15]), .QB (
         \$dummy [217]), .D (nx19573), .CLK (clk), .R (rst)) ;
    latch lat_label_10_input_15 (.Q (label_10_input_15), .D (nx9428), .CLK (
          nx34519)) ;
    dffr reg_label_10_input_state_machine_15 (.Q (
         label_10_input_state_machine_15), .QB (\$dummy [218]), .D (nx19563), .CLK (
         clk), .R (rst)) ;
    xnor2 ix9425 (.Y (nx9424), .A0 (nx9420), .A1 (nx28150)) ;
    oai22 ix9421 (.Y (nx9420), .A0 (nx27586), .A1 (nx27758), .B0 (nx27760), .B1 (
          nx27554)) ;
    oai21 ix19614 (.Y (nx19613), .A0 (nx28155), .A1 (nx34763), .B0 (nx28157)) ;
    dff max_calc_reg_comparator_fifth_inp1_15 (.Q (\$dummy [219]), .QB (nx28155)
        , .D (nx19613), .CLK (clk)) ;
    nand03 ix28158 (.Y (nx28157), .A0 (label_9_output[15]), .A1 (nx34745), .A2 (
           nx34765)) ;
    dffr labelsregfile_label9_loop1_15_fx_reg_q (.Q (label_9_output[15]), .QB (
         \$dummy [220]), .D (nx19603), .CLK (clk), .R (rst)) ;
    latch lat_label_9_input_15 (.Q (label_9_input_15), .D (nx9468), .CLK (
          nx34519)) ;
    dffr reg_label_9_input_state_machine_15 (.Q (label_9_input_state_machine_15)
         , .QB (\$dummy [221]), .D (nx19593), .CLK (clk), .R (rst)) ;
    xnor2 ix9465 (.Y (nx9464), .A0 (nx9460), .A1 (nx28168)) ;
    oai22 ix9461 (.Y (nx9460), .A0 (nx27775), .A1 (nx27947), .B0 (nx27949), .B1 (
          nx27115)) ;
    dff max_calc_reg_comparator_first_inp2_0 (.Q (
        max_calc_comparator_first_inp2_0), .QB (nx33288), .D (nx25473), .CLK (
        clk)) ;
    dffr labelsregfile_label2_loop1_0_fx_reg_q (.Q (label_2_output[0]), .QB (
         \$dummy [222]), .D (nx16373), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_0 (.Q (label_2_input_0), .D (nx4420), .CLK (nx34519)
          ) ;
    oai21 ix4421 (.Y (nx4420), .A0 (nx28183), .A1 (nx34419), .B0 (nx28187)) ;
    dffr reg_label_2_input_state_machine_0 (.Q (label_2_input_state_machine_0), 
         .QB (nx28183), .D (nx16363), .CLK (clk), .R (rst)) ;
    oai21 ix28188 (.Y (nx28187), .A0 (nx35727), .A1 (label_2_output[0]), .B0 (
          nx4408)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_1_1), .QB (\$dummy [223]), .D (nx16343)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_1_2), .QB (nx28608), .D (nx16333), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_1_3), .QB (\$dummy [224]), .D (nx16323)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_1_4), .QB (nx28606), .D (nx16313), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_1_5), .QB (\$dummy [225]), .D (nx16303)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_1_6), .QB (nx28604), .D (nx16293), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_1_7), .QB (\$dummy [226]), .D (nx16283)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_1_8), .QB (nx28602), .D (nx16273), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_1_9), .QB (\$dummy [227]), .D (nx16263)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_1_10), .QB (nx28600), .D (nx16253), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_1_11), .QB (\$dummy [228]), .D (nx16243)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_1_12), .QB (nx28598), .D (nx16233), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_1_13), .QB (\$dummy [229]), .D (nx16223)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_1_14), .QB (nx28596), .D (nx16213), .CLK (
         clk), .R (rst)) ;
    aoi22 ix28237 (.Y (nx28236), .A0 (mdr_data_out[15]), .A1 (nx34635), .B0 (
          nx4206), .B1 (nx4212)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_reg_output_0), .QB (\$dummy [230]), .D (
         nx15853), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_1_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_1_shift_Reg_count_0), .QB (\$dummy [231]), .D (
            nx15839), .CLK (clk), .S (nx34475)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_reg_output_9), .QB (\$dummy [232]), .D (
         nx16033), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_9), .QB (\$dummy [233]), .D (
         nx16023), .CLK (clk), .R (nx34473)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_8), .QB (\$dummy [234]), .D (
         nx16013), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_8), .QB (\$dummy [235]), .D (
         nx16003), .CLK (clk), .R (nx34473)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_7), .QB (\$dummy [236]), .D (
         nx15993), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_7), .QB (\$dummy [237]), .D (
         nx15983), .CLK (clk), .R (nx34473)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_6), .QB (\$dummy [238]), .D (
         nx15973), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_6), .QB (\$dummy [239]), .D (
         nx15963), .CLK (clk), .R (nx34473)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_5), .QB (\$dummy [240]), .D (
         nx15953), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_5), .QB (\$dummy [241]), .D (
         nx15943), .CLK (clk), .R (nx34473)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_4), .QB (\$dummy [242]), .D (
         nx15933), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_4), .QB (\$dummy [243]), .D (
         nx15923), .CLK (clk), .R (nx34473)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_3), .QB (\$dummy [244]), .D (
         nx15913), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_3), .QB (\$dummy [245]), .D (
         nx15903), .CLK (clk), .R (nx34473)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_2), .QB (\$dummy [246]), .D (
         nx15893), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_2), .QB (\$dummy [247]), .D (
         nx15883), .CLK (clk), .R (nx34471)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_1_shift_Reg_output_1), .QB (\$dummy [248]), .D (
         nx15873), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_1_shift_Reg_count_1), .QB (\$dummy [249]), .D (
         nx15863), .CLK (clk), .R (nx34471)) ;
    nand02 ix15834 (.Y (nx15833), .A0 (nx35815), .A1 (nx34621)) ;
    dffs_ni booth_booth_integrtaion_1_shift_Reg_reg_en (.Q (\$dummy [250]), .QB (
            nx28283), .D (nx15833), .CLK (clk), .S (nx34471)) ;
    nand02 ix4207 (.Y (nx4206), .A0 (nx28304), .A1 (nx28316)) ;
    oai21 ix28305 (.Y (nx28304), .A0 (nx34649), .A1 (nx34643), .B0 (
          mdr_data_out[32])) ;
    oai21 ix16044 (.Y (nx16043), .A0 (nx28309), .A1 (nx35373), .B0 (nx28311)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [251]), .QB (
         nx28309), .D (nx16043), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [252]), .QB (
         nx28313), .D (nx16353), .CLK (clk), .R (rst)) ;
    xnor2 ix28321 (.Y (nx28320), .A0 (nx3676), .A1 (nx13017)) ;
    oai21 ix16184 (.Y (nx16183), .A0 (nx28326), .A1 (nx35373), .B0 (nx28328)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_17), .QB (nx28326), .D (nx16183)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28329 (.Y (nx28328), .A0 (nx35381), .A1 (nx4184), .A2 (nx36077)) ;
    xnor2 ix4185 (.Y (nx4184), .A0 (nx28331), .A1 (nx13018)) ;
    aoi22 ix28332 (.Y (nx28331), .A0 (booth_booth_integrtaion_1_booth_output_17)
          , .A1 (nx3700), .B0 (nx3676), .B1 (nx13017)) ;
    nand02 ix3685 (.Y (nx3684), .A0 (mdr_data_out[33]), .A1 (mdr_data_out[32])
           ) ;
    or02 ix28336 (.Y (nx28335), .A0 (mdr_data_out[32]), .A1 (mdr_data_out[33])
         ) ;
    xnor2 ix28342 (.Y (nx28341), .A0 (nx3728), .A1 (nx13019)) ;
    oai22 ix3729 (.Y (nx3728), .A0 (nx28331), .A1 (nx28344), .B0 (nx28351), .B1 (
          nx35385)) ;
    aoi32 ix28347 (.Y (nx28346), .A0 (nx3710), .A1 (nx34649), .A2 (nx28349), .B0 (
          mdr_data_out[34]), .B1 (nx34643)) ;
    oai21 ix3711 (.Y (nx3710), .A0 (mdr_data_out[32]), .A1 (mdr_data_out[33]), .B0 (
          mdr_data_out[34])) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_18), .QB (nx28351), .D (nx16173)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16164 (.Y (nx16163), .A0 (nx28356), .A1 (nx35373), .B0 (nx28358)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_19), .QB (nx28356), .D (nx16163)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28359 (.Y (nx28358), .A0 (nx35381), .A1 (nx4160), .A2 (nx36077)) ;
    xnor2 ix4161 (.Y (nx4160), .A0 (nx28361), .A1 (nx13021)) ;
    aoi22 ix28362 (.Y (nx28361), .A0 (booth_booth_integrtaion_1_booth_output_19)
          , .A1 (nx3748), .B0 (nx3728), .B1 (nx13019)) ;
    nor02ii ix28365 (.Y (nx28364), .A0 (nx3714), .A1 (mdr_data_out[35])) ;
    nor03_2x ix3715 (.Y (nx3714), .A0 (mdr_data_out[34]), .A1 (mdr_data_out[32])
             , .A2 (mdr_data_out[33])) ;
    nor04 ix3739 (.Y (nx3738), .A0 (mdr_data_out[35]), .A1 (mdr_data_out[34]), .A2 (
          mdr_data_out[32]), .A3 (mdr_data_out[33])) ;
    xnor2 ix28379 (.Y (nx28378), .A0 (nx3776), .A1 (nx13023)) ;
    oai22 ix3777 (.Y (nx3776), .A0 (nx28361), .A1 (nx28381), .B0 (nx28390), .B1 (
          nx35387)) ;
    aoi32 ix28384 (.Y (nx28383), .A0 (nx3758), .A1 (nx34649), .A2 (nx28388), .B0 (
          mdr_data_out[36]), .B1 (nx34643)) ;
    nand02 ix3759 (.Y (nx3758), .A0 (nx28386), .A1 (mdr_data_out[36])) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_20), .QB (nx28390), .D (nx16153)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16144 (.Y (nx16143), .A0 (nx28395), .A1 (nx35373), .B0 (nx28397)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_21), .QB (nx28395), .D (nx16143)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28398 (.Y (nx28397), .A0 (nx35381), .A1 (nx4136), .A2 (nx36077)) ;
    xnor2 ix4137 (.Y (nx4136), .A0 (nx28400), .A1 (nx13025)) ;
    aoi22 ix28401 (.Y (nx28400), .A0 (booth_booth_integrtaion_1_booth_output_21)
          , .A1 (nx3796), .B0 (nx3776), .B1 (nx13023)) ;
    nor02ii ix28404 (.Y (nx28403), .A0 (nx3762), .A1 (mdr_data_out[37])) ;
    nor02ii ix3763 (.Y (nx3762), .A0 (mdr_data_out[36]), .A1 (nx3738)) ;
    nor02ii ix3787 (.Y (nx3786), .A0 (mdr_data_out[37]), .A1 (nx3762)) ;
    xnor2 ix28414 (.Y (nx28413), .A0 (nx3824), .A1 (nx13026)) ;
    oai22 ix3825 (.Y (nx3824), .A0 (nx28400), .A1 (nx28416), .B0 (nx28425), .B1 (
          nx35389)) ;
    aoi32 ix28419 (.Y (nx28418), .A0 (nx3806), .A1 (nx34649), .A2 (nx28423), .B0 (
          mdr_data_out[38]), .B1 (nx34643)) ;
    nand02 ix3807 (.Y (nx3806), .A0 (nx28421), .A1 (mdr_data_out[38])) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_22), .QB (nx28425), .D (nx16133)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16124 (.Y (nx16123), .A0 (nx28430), .A1 (nx35373), .B0 (nx28432)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_23), .QB (nx28430), .D (nx16123)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28433 (.Y (nx28432), .A0 (nx35381), .A1 (nx4112), .A2 (nx35375)) ;
    xnor2 ix4113 (.Y (nx4112), .A0 (nx28435), .A1 (nx13027)) ;
    aoi22 ix28436 (.Y (nx28435), .A0 (booth_booth_integrtaion_1_booth_output_23)
          , .A1 (nx3844), .B0 (nx3824), .B1 (nx13026)) ;
    nor02ii ix28439 (.Y (nx28438), .A0 (nx3810), .A1 (mdr_data_out[39])) ;
    nor02ii ix3811 (.Y (nx3810), .A0 (mdr_data_out[38]), .A1 (nx3786)) ;
    nor02ii ix3835 (.Y (nx3834), .A0 (mdr_data_out[39]), .A1 (nx3810)) ;
    xnor2 ix28449 (.Y (nx28448), .A0 (nx3872), .A1 (nx13029)) ;
    oai22 ix3873 (.Y (nx3872), .A0 (nx28435), .A1 (nx28451), .B0 (nx28460), .B1 (
          nx35391)) ;
    aoi32 ix28454 (.Y (nx28453), .A0 (nx3854), .A1 (nx34649), .A2 (nx28458), .B0 (
          mdr_data_out[40]), .B1 (nx34643)) ;
    nand02 ix3855 (.Y (nx3854), .A0 (nx28456), .A1 (mdr_data_out[40])) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_24), .QB (nx28460), .D (nx16113)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16104 (.Y (nx16103), .A0 (nx28465), .A1 (nx35375), .B0 (nx28467)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_25), .QB (nx28465), .D (nx16103)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28468 (.Y (nx28467), .A0 (nx35381), .A1 (nx4088), .A2 (nx35375)) ;
    xnor2 ix4089 (.Y (nx4088), .A0 (nx28470), .A1 (nx13031)) ;
    aoi22 ix28471 (.Y (nx28470), .A0 (booth_booth_integrtaion_1_booth_output_25)
          , .A1 (nx3892), .B0 (nx3872), .B1 (nx13029)) ;
    nor02ii ix28474 (.Y (nx28473), .A0 (nx3858), .A1 (mdr_data_out[41])) ;
    nor02ii ix3859 (.Y (nx3858), .A0 (mdr_data_out[40]), .A1 (nx3834)) ;
    nor02ii ix3883 (.Y (nx3882), .A0 (mdr_data_out[41]), .A1 (nx3858)) ;
    xnor2 ix28484 (.Y (nx28483), .A0 (nx3920), .A1 (nx13033)) ;
    oai22 ix3921 (.Y (nx3920), .A0 (nx28470), .A1 (nx28486), .B0 (nx28495), .B1 (
          nx35393)) ;
    aoi32 ix28489 (.Y (nx28488), .A0 (nx3902), .A1 (nx34649), .A2 (nx28493), .B0 (
          mdr_data_out[42]), .B1 (nx34643)) ;
    nand02 ix3903 (.Y (nx3902), .A0 (nx28491), .A1 (mdr_data_out[42])) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_26), .QB (nx28495), .D (nx16093)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16084 (.Y (nx16083), .A0 (nx28500), .A1 (nx35375), .B0 (nx28502)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_27), .QB (nx28500), .D (nx16083)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28503 (.Y (nx28502), .A0 (nx35381), .A1 (nx4064), .A2 (nx35375)) ;
    xnor2 ix4065 (.Y (nx4064), .A0 (nx28505), .A1 (nx13035)) ;
    aoi22 ix28506 (.Y (nx28505), .A0 (booth_booth_integrtaion_1_booth_output_27)
          , .A1 (nx3940), .B0 (nx3920), .B1 (nx13033)) ;
    nor02ii ix28509 (.Y (nx28508), .A0 (nx3906), .A1 (mdr_data_out[43])) ;
    nor02ii ix3907 (.Y (nx3906), .A0 (mdr_data_out[42]), .A1 (nx3882)) ;
    nor02ii ix3931 (.Y (nx3930), .A0 (mdr_data_out[43]), .A1 (nx3906)) ;
    xnor2 ix28519 (.Y (nx28518), .A0 (nx3968), .A1 (nx13037)) ;
    oai22 ix3969 (.Y (nx3968), .A0 (nx28505), .A1 (nx28521), .B0 (nx28530), .B1 (
          nx35395)) ;
    aoi32 ix28524 (.Y (nx28523), .A0 (nx3950), .A1 (nx34649), .A2 (nx28528), .B0 (
          mdr_data_out[44]), .B1 (nx34643)) ;
    nand02 ix3951 (.Y (nx3950), .A0 (nx28526), .A1 (mdr_data_out[44])) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_28), .QB (nx28530), .D (nx16073)
         , .CLK (clk), .R (rst)) ;
    oai21 ix16064 (.Y (nx16063), .A0 (nx28535), .A1 (nx35375), .B0 (nx28537)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_29), .QB (nx28535), .D (nx16063)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28538 (.Y (nx28537), .A0 (nx36085), .A1 (nx4040), .A2 (nx35375)) ;
    xnor2 ix4041 (.Y (nx4040), .A0 (nx28540), .A1 (nx13039)) ;
    aoi22 ix28541 (.Y (nx28540), .A0 (booth_booth_integrtaion_1_booth_output_29)
          , .A1 (nx3988), .B0 (nx3968), .B1 (nx13037)) ;
    nor02ii ix28544 (.Y (nx28543), .A0 (nx3954), .A1 (mdr_data_out[45])) ;
    nor02ii ix3955 (.Y (nx3954), .A0 (mdr_data_out[44]), .A1 (nx3930)) ;
    nor02ii ix3979 (.Y (nx3978), .A0 (mdr_data_out[45]), .A1 (nx3954)) ;
    xnor2 ix28554 (.Y (nx28553), .A0 (nx4016), .A1 (nx4026)) ;
    oai22 ix4017 (.Y (nx4016), .A0 (nx28540), .A1 (nx28556), .B0 (nx28565), .B1 (
          nx35397)) ;
    aoi32 ix28559 (.Y (nx28558), .A0 (nx3998), .A1 (nx34651), .A2 (nx28563), .B0 (
          mdr_data_out[46]), .B1 (nx34645)) ;
    nand02 ix3999 (.Y (nx3998), .A0 (nx28561), .A1 (mdr_data_out[46])) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_31), .QB (nx28565), .D (nx16053)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix28569 (.Y (nx28568), .A0 (mdr_data_out[47]), .A1 (nx34645), .B0 (
          nx34651), .B1 (nx4018)) ;
    xnor2 ix4019 (.Y (nx4018), .A0 (mdr_data_out[47]), .A1 (nx4002)) ;
    nor02ii ix4003 (.Y (nx4002), .A0 (mdr_data_out[46]), .A1 (nx3978)) ;
    aoi32 ix28573 (.Y (nx28572), .A0 (nx3974), .A1 (nx34651), .A2 (nx28561), .B0 (
          mdr_data_out[45]), .B1 (nx34645)) ;
    aoi32 ix28576 (.Y (nx28575), .A0 (nx3926), .A1 (nx34651), .A2 (nx28526), .B0 (
          mdr_data_out[43]), .B1 (nx34645)) ;
    aoi32 ix28579 (.Y (nx28578), .A0 (nx3878), .A1 (nx34651), .A2 (nx28491), .B0 (
          mdr_data_out[41]), .B1 (nx34645)) ;
    aoi32 ix28582 (.Y (nx28581), .A0 (nx3830), .A1 (nx34651), .A2 (nx28456), .B0 (
          mdr_data_out[39]), .B1 (nx34645)) ;
    aoi32 ix28585 (.Y (nx28584), .A0 (nx3782), .A1 (nx34651), .A2 (nx28421), .B0 (
          mdr_data_out[37]), .B1 (nx34645)) ;
    aoi32 ix28588 (.Y (nx28587), .A0 (nx3734), .A1 (nx3670), .A2 (nx28386), .B0 (
          mdr_data_out[35]), .B1 (nx34647)) ;
    aoi32 ix28591 (.Y (nx28590), .A0 (nx3684), .A1 (nx3670), .A2 (nx28335), .B0 (
          mdr_data_out[33]), .B1 (nx34647)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_1_booth_output_16), .QB (nx28316), .D (nx16193)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_1_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_1_15), .QB (nx28594), .D (nx16203), .CLK (
         clk), .R (rst)) ;
    aoi21 ix4409 (.Y (nx4408), .A0 (label_2_output[0]), .A1 (nx35727), .B0 (
          nx36387)) ;
    dff max_calc_reg_ans2_0 (.Q (max_calc_ans2_0), .QB (\$dummy [253]), .D (
        nx25443), .CLK (clk)) ;
    oai21 ix24274 (.Y (nx24273), .A0 (nx28617), .A1 (nx34765), .B0 (nx28619)) ;
    dff max_calc_reg_comparator_second_inp1_0 (.Q (
        max_calc_comparator_second_inp1_0), .QB (nx28617), .D (nx24273), .CLK (
        clk)) ;
    nand03 ix28620 (.Y (nx28619), .A0 (nx36389), .A1 (nx16932), .A2 (nx34783)) ;
    dffr labelsregfile_label3_loop1_0_fx_reg_q (.Q (label_3_output[0]), .QB (
         \$dummy [254]), .D (nx15523), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_0 (.Q (label_3_input_0), .D (nx3082), .CLK (nx34519)
          ) ;
    oai21 ix3083 (.Y (nx3082), .A0 (nx28626), .A1 (nx34419), .B0 (nx28630)) ;
    dffr reg_label_3_input_state_machine_0 (.Q (label_3_input_state_machine_0), 
         .QB (nx28626), .D (nx15513), .CLK (clk), .R (rst)) ;
    oai21 ix28631 (.Y (nx28630), .A0 (nx35723), .A1 (label_3_output[0]), .B0 (
          nx3070)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_2_1), .QB (\$dummy [255]), .D (nx15493)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_2_2), .QB (nx29051), .D (nx15483), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_2_3), .QB (\$dummy [256]), .D (nx15473)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_2_4), .QB (nx29049), .D (nx15463), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_2_5), .QB (\$dummy [257]), .D (nx15453)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_2_6), .QB (nx29047), .D (nx15443), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_2_7), .QB (\$dummy [258]), .D (nx15433)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_2_8), .QB (nx29045), .D (nx15423), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_2_9), .QB (\$dummy [259]), .D (nx15413)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_2_10), .QB (nx29043), .D (nx15403), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_2_11), .QB (\$dummy [260]), .D (nx15393)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_2_12), .QB (nx29041), .D (nx15383), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_2_13), .QB (\$dummy [261]), .D (nx15373)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_2_14), .QB (nx29039), .D (nx15363), .CLK (
         clk), .R (rst)) ;
    aoi22 ix28680 (.Y (nx28679), .A0 (mdr_data_out[15]), .A1 (nx34603), .B0 (
          nx2868), .B1 (nx2874)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_reg_output_0), .QB (\$dummy [262]), .D (
         nx15003), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_2_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_2_shift_Reg_count_0), .QB (\$dummy [263]), .D (
            nx14989), .CLK (clk), .S (nx34477)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_reg_output_9), .QB (\$dummy [264]), .D (
         nx15183), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_9), .QB (\$dummy [265]), .D (
         nx15173), .CLK (clk), .R (nx34477)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_8), .QB (\$dummy [266]), .D (
         nx15163), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_8), .QB (\$dummy [267]), .D (
         nx15153), .CLK (clk), .R (nx34477)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_7), .QB (\$dummy [268]), .D (
         nx15143), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_7), .QB (\$dummy [269]), .D (
         nx15133), .CLK (clk), .R (nx34477)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_6), .QB (\$dummy [270]), .D (
         nx15123), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_6), .QB (\$dummy [271]), .D (
         nx15113), .CLK (clk), .R (nx34477)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_5), .QB (\$dummy [272]), .D (
         nx15103), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_5), .QB (\$dummy [273]), .D (
         nx15093), .CLK (clk), .R (nx34475)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_4), .QB (\$dummy [274]), .D (
         nx15083), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_4), .QB (\$dummy [275]), .D (
         nx15073), .CLK (clk), .R (nx34475)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_3), .QB (\$dummy [276]), .D (
         nx15063), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_3), .QB (\$dummy [277]), .D (
         nx15053), .CLK (clk), .R (nx34475)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_2), .QB (\$dummy [278]), .D (
         nx15043), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_2), .QB (\$dummy [279]), .D (
         nx15033), .CLK (clk), .R (nx34475)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_2_shift_Reg_output_1), .QB (\$dummy [280]), .D (
         nx15023), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_2_shift_Reg_count_1), .QB (\$dummy [281]), .D (
         nx15013), .CLK (clk), .R (nx34475)) ;
    nand02 ix14984 (.Y (nx14983), .A0 (nx35819), .A1 (nx34589)) ;
    dffs_ni booth_booth_integrtaion_2_shift_Reg_reg_en (.Q (\$dummy [282]), .QB (
            nx28726), .D (nx14983), .CLK (clk), .S (nx34475)) ;
    nand02 ix2869 (.Y (nx2868), .A0 (nx28747), .A1 (nx28759)) ;
    oai21 ix28748 (.Y (nx28747), .A0 (nx34617), .A1 (nx34611), .B0 (
          mdr_data_out[48])) ;
    oai21 ix15194 (.Y (nx15193), .A0 (nx28752), .A1 (nx35399), .B0 (nx28754)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [283]), .QB (
         nx28752), .D (nx15193), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [284]), .QB (
         nx28756), .D (nx15503), .CLK (clk), .R (rst)) ;
    xnor2 ix28764 (.Y (nx28763), .A0 (nx2338), .A1 (nx12965)) ;
    oai21 ix15334 (.Y (nx15333), .A0 (nx28769), .A1 (nx35399), .B0 (nx28771)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_17), .QB (nx28769), .D (nx15333)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28772 (.Y (nx28771), .A0 (nx35407), .A1 (nx2846), .A2 (nx36093)) ;
    xnor2 ix2847 (.Y (nx2846), .A0 (nx28774), .A1 (nx12967)) ;
    aoi22 ix28775 (.Y (nx28774), .A0 (booth_booth_integrtaion_2_booth_output_17)
          , .A1 (nx2362), .B0 (nx2338), .B1 (nx12965)) ;
    nand02 ix2347 (.Y (nx2346), .A0 (mdr_data_out[49]), .A1 (mdr_data_out[48])
           ) ;
    or02 ix28779 (.Y (nx28778), .A0 (mdr_data_out[48]), .A1 (mdr_data_out[49])
         ) ;
    xnor2 ix28785 (.Y (nx28784), .A0 (nx2390), .A1 (nx12969)) ;
    oai22 ix2391 (.Y (nx2390), .A0 (nx28774), .A1 (nx28787), .B0 (nx28794), .B1 (
          nx35411)) ;
    aoi32 ix28790 (.Y (nx28789), .A0 (nx2372), .A1 (nx34617), .A2 (nx28792), .B0 (
          mdr_data_out[50]), .B1 (nx34611)) ;
    oai21 ix2373 (.Y (nx2372), .A0 (mdr_data_out[48]), .A1 (mdr_data_out[49]), .B0 (
          mdr_data_out[50])) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_18), .QB (nx28794), .D (nx15323)
         , .CLK (clk), .R (rst)) ;
    oai21 ix15314 (.Y (nx15313), .A0 (nx28799), .A1 (nx35399), .B0 (nx28801)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_19), .QB (nx28799), .D (nx15313)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28802 (.Y (nx28801), .A0 (nx35407), .A1 (nx2822), .A2 (nx36093)) ;
    xnor2 ix2823 (.Y (nx2822), .A0 (nx28804), .A1 (nx12970)) ;
    aoi22 ix28805 (.Y (nx28804), .A0 (booth_booth_integrtaion_2_booth_output_19)
          , .A1 (nx2410), .B0 (nx2390), .B1 (nx12969)) ;
    nor02ii ix28808 (.Y (nx28807), .A0 (nx2376), .A1 (mdr_data_out[51])) ;
    nor03_2x ix2377 (.Y (nx2376), .A0 (mdr_data_out[50]), .A1 (mdr_data_out[48])
             , .A2 (mdr_data_out[49])) ;
    nor04 ix2401 (.Y (nx2400), .A0 (mdr_data_out[51]), .A1 (mdr_data_out[50]), .A2 (
          mdr_data_out[48]), .A3 (mdr_data_out[49])) ;
    xnor2 ix28822 (.Y (nx28821), .A0 (nx2438), .A1 (nx12971)) ;
    oai22 ix2439 (.Y (nx2438), .A0 (nx28804), .A1 (nx28824), .B0 (nx28833), .B1 (
          nx35413)) ;
    aoi32 ix28827 (.Y (nx28826), .A0 (nx2420), .A1 (nx34617), .A2 (nx28831), .B0 (
          mdr_data_out[52]), .B1 (nx34611)) ;
    nand02 ix2421 (.Y (nx2420), .A0 (nx28829), .A1 (mdr_data_out[52])) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_20), .QB (nx28833), .D (nx15303)
         , .CLK (clk), .R (rst)) ;
    oai21 ix15294 (.Y (nx15293), .A0 (nx28838), .A1 (nx35399), .B0 (nx28840)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_21), .QB (nx28838), .D (nx15293)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28841 (.Y (nx28840), .A0 (nx35407), .A1 (nx2798), .A2 (nx36093)) ;
    xnor2 ix2799 (.Y (nx2798), .A0 (nx28843), .A1 (nx12973)) ;
    aoi22 ix28844 (.Y (nx28843), .A0 (booth_booth_integrtaion_2_booth_output_21)
          , .A1 (nx2458), .B0 (nx2438), .B1 (nx12971)) ;
    nor02ii ix28847 (.Y (nx28846), .A0 (nx2424), .A1 (mdr_data_out[53])) ;
    nor02ii ix2425 (.Y (nx2424), .A0 (mdr_data_out[52]), .A1 (nx2400)) ;
    nor02ii ix2449 (.Y (nx2448), .A0 (mdr_data_out[53]), .A1 (nx2424)) ;
    xnor2 ix28857 (.Y (nx28856), .A0 (nx2486), .A1 (nx12975)) ;
    oai22 ix2487 (.Y (nx2486), .A0 (nx28843), .A1 (nx28859), .B0 (nx28868), .B1 (
          nx35415)) ;
    aoi32 ix28862 (.Y (nx28861), .A0 (nx2468), .A1 (nx34617), .A2 (nx28866), .B0 (
          mdr_data_out[54]), .B1 (nx34611)) ;
    nand02 ix2469 (.Y (nx2468), .A0 (nx28864), .A1 (mdr_data_out[54])) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_22), .QB (nx28868), .D (nx15283)
         , .CLK (clk), .R (rst)) ;
    oai21 ix15274 (.Y (nx15273), .A0 (nx28873), .A1 (nx35399), .B0 (nx28875)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_23), .QB (nx28873), .D (nx15273)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28876 (.Y (nx28875), .A0 (nx35407), .A1 (nx2774), .A2 (nx35401)) ;
    xnor2 ix2775 (.Y (nx2774), .A0 (nx28878), .A1 (nx12977)) ;
    aoi22 ix28879 (.Y (nx28878), .A0 (booth_booth_integrtaion_2_booth_output_23)
          , .A1 (nx2506), .B0 (nx2486), .B1 (nx12975)) ;
    nor02ii ix28882 (.Y (nx28881), .A0 (nx2472), .A1 (mdr_data_out[55])) ;
    nor02ii ix2473 (.Y (nx2472), .A0 (mdr_data_out[54]), .A1 (nx2448)) ;
    nor02ii ix2497 (.Y (nx2496), .A0 (mdr_data_out[55]), .A1 (nx2472)) ;
    xnor2 ix28892 (.Y (nx28891), .A0 (nx2534), .A1 (nx12978)) ;
    oai22 ix2535 (.Y (nx2534), .A0 (nx28878), .A1 (nx28894), .B0 (nx28903), .B1 (
          nx35417)) ;
    aoi32 ix28897 (.Y (nx28896), .A0 (nx2516), .A1 (nx34617), .A2 (nx28901), .B0 (
          mdr_data_out[56]), .B1 (nx34611)) ;
    nand02 ix2517 (.Y (nx2516), .A0 (nx28899), .A1 (mdr_data_out[56])) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_24), .QB (nx28903), .D (nx15263)
         , .CLK (clk), .R (rst)) ;
    oai21 ix15254 (.Y (nx15253), .A0 (nx28908), .A1 (nx35401), .B0 (nx28910)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_25), .QB (nx28908), .D (nx15253)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28911 (.Y (nx28910), .A0 (nx35407), .A1 (nx2750), .A2 (nx35401)) ;
    xnor2 ix2751 (.Y (nx2750), .A0 (nx28913), .A1 (nx12979)) ;
    aoi22 ix28914 (.Y (nx28913), .A0 (booth_booth_integrtaion_2_booth_output_25)
          , .A1 (nx2554), .B0 (nx2534), .B1 (nx12978)) ;
    nor02ii ix28917 (.Y (nx28916), .A0 (nx2520), .A1 (mdr_data_out[57])) ;
    nor02ii ix2521 (.Y (nx2520), .A0 (mdr_data_out[56]), .A1 (nx2496)) ;
    nor02ii ix2545 (.Y (nx2544), .A0 (mdr_data_out[57]), .A1 (nx2520)) ;
    xnor2 ix28927 (.Y (nx28926), .A0 (nx2582), .A1 (nx12981)) ;
    oai22 ix2583 (.Y (nx2582), .A0 (nx28913), .A1 (nx28929), .B0 (nx28938), .B1 (
          nx35419)) ;
    aoi32 ix28932 (.Y (nx28931), .A0 (nx2564), .A1 (nx34617), .A2 (nx28936), .B0 (
          mdr_data_out[58]), .B1 (nx34611)) ;
    nand02 ix2565 (.Y (nx2564), .A0 (nx28934), .A1 (mdr_data_out[58])) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_26), .QB (nx28938), .D (nx15243)
         , .CLK (clk), .R (rst)) ;
    oai21 ix15234 (.Y (nx15233), .A0 (nx28943), .A1 (nx35401), .B0 (nx28945)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_27), .QB (nx28943), .D (nx15233)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28946 (.Y (nx28945), .A0 (nx35407), .A1 (nx2726), .A2 (nx35401)) ;
    xnor2 ix2727 (.Y (nx2726), .A0 (nx28948), .A1 (nx12983)) ;
    aoi22 ix28949 (.Y (nx28948), .A0 (booth_booth_integrtaion_2_booth_output_27)
          , .A1 (nx2602), .B0 (nx2582), .B1 (nx12981)) ;
    nor02ii ix28952 (.Y (nx28951), .A0 (nx2568), .A1 (mdr_data_out[59])) ;
    nor02ii ix2569 (.Y (nx2568), .A0 (mdr_data_out[58]), .A1 (nx2544)) ;
    nor02ii ix2593 (.Y (nx2592), .A0 (mdr_data_out[59]), .A1 (nx2568)) ;
    xnor2 ix28962 (.Y (nx28961), .A0 (nx2630), .A1 (nx12985)) ;
    oai22 ix2631 (.Y (nx2630), .A0 (nx28948), .A1 (nx28964), .B0 (nx28973), .B1 (
          nx35421)) ;
    aoi32 ix28967 (.Y (nx28966), .A0 (nx2612), .A1 (nx34617), .A2 (nx28971), .B0 (
          mdr_data_out[60]), .B1 (nx34611)) ;
    nand02 ix2613 (.Y (nx2612), .A0 (nx28969), .A1 (mdr_data_out[60])) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_28), .QB (nx28973), .D (nx15223)
         , .CLK (clk), .R (rst)) ;
    oai21 ix15214 (.Y (nx15213), .A0 (nx28978), .A1 (nx35401), .B0 (nx28980)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_29), .QB (nx28978), .D (nx15213)
         , .CLK (clk), .R (rst)) ;
    nand03 ix28981 (.Y (nx28980), .A0 (nx36101), .A1 (nx2702), .A2 (nx35401)) ;
    xnor2 ix2703 (.Y (nx2702), .A0 (nx28983), .A1 (nx12987)) ;
    aoi22 ix28984 (.Y (nx28983), .A0 (booth_booth_integrtaion_2_booth_output_29)
          , .A1 (nx2650), .B0 (nx2630), .B1 (nx12985)) ;
    nor02ii ix28987 (.Y (nx28986), .A0 (nx2616), .A1 (mdr_data_out[61])) ;
    nor02ii ix2617 (.Y (nx2616), .A0 (mdr_data_out[60]), .A1 (nx2592)) ;
    nor02ii ix2641 (.Y (nx2640), .A0 (mdr_data_out[61]), .A1 (nx2616)) ;
    xnor2 ix28997 (.Y (nx28996), .A0 (nx2678), .A1 (nx2688)) ;
    oai22 ix2679 (.Y (nx2678), .A0 (nx28983), .A1 (nx28999), .B0 (nx29008), .B1 (
          nx35423)) ;
    aoi32 ix29002 (.Y (nx29001), .A0 (nx2660), .A1 (nx34619), .A2 (nx29006), .B0 (
          mdr_data_out[62]), .B1 (nx34613)) ;
    nand02 ix2661 (.Y (nx2660), .A0 (nx29004), .A1 (mdr_data_out[62])) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_31), .QB (nx29008), .D (nx15203)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix29012 (.Y (nx29011), .A0 (mdr_data_out[63]), .A1 (nx34613), .B0 (
          nx34619), .B1 (nx2680)) ;
    xnor2 ix2681 (.Y (nx2680), .A0 (mdr_data_out[63]), .A1 (nx2664)) ;
    nor02ii ix2665 (.Y (nx2664), .A0 (mdr_data_out[62]), .A1 (nx2640)) ;
    aoi32 ix29016 (.Y (nx29015), .A0 (nx2636), .A1 (nx34619), .A2 (nx29004), .B0 (
          mdr_data_out[61]), .B1 (nx34613)) ;
    aoi32 ix29019 (.Y (nx29018), .A0 (nx2588), .A1 (nx34619), .A2 (nx28969), .B0 (
          mdr_data_out[59]), .B1 (nx34613)) ;
    aoi32 ix29022 (.Y (nx29021), .A0 (nx2540), .A1 (nx34619), .A2 (nx28934), .B0 (
          mdr_data_out[57]), .B1 (nx34613)) ;
    aoi32 ix29025 (.Y (nx29024), .A0 (nx2492), .A1 (nx34619), .A2 (nx28899), .B0 (
          mdr_data_out[55]), .B1 (nx34613)) ;
    aoi32 ix29028 (.Y (nx29027), .A0 (nx2444), .A1 (nx34619), .A2 (nx28864), .B0 (
          mdr_data_out[53]), .B1 (nx34613)) ;
    aoi32 ix29031 (.Y (nx29030), .A0 (nx2396), .A1 (nx2332), .A2 (nx28829), .B0 (
          mdr_data_out[51]), .B1 (nx34615)) ;
    aoi32 ix29034 (.Y (nx29033), .A0 (nx2346), .A1 (nx2332), .A2 (nx28778), .B0 (
          mdr_data_out[49]), .B1 (nx34615)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_2_booth_output_16), .QB (nx28759), .D (nx15343)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_2_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_2_15), .QB (nx29037), .D (nx15353), .CLK (
         clk), .R (rst)) ;
    aoi21 ix3071 (.Y (nx3070), .A0 (label_3_output[0]), .A1 (nx35723), .B0 (
          nx36387)) ;
    oai21 ix21594 (.Y (nx21593), .A0 (nx29061), .A1 (nx34765), .B0 (nx29063)) ;
    dff max_calc_reg_comparator_third_inp1_0 (.Q (
        max_calc_comparator_third_inp1_0), .QB (nx29061), .D (nx21593), .CLK (
        clk)) ;
    nand03 ix29064 (.Y (nx29063), .A0 (label_5_output[0]), .A1 (nx35453), .A2 (
           nx34765)) ;
    dffr labelsregfile_label5_loop1_0_fx_reg_q (.Q (label_5_output[0]), .QB (
         \$dummy [285]), .D (nx20193), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_0 (.Q (label_5_input_0), .D (nx10396), .CLK (nx34521
          )) ;
    oai21 ix10397 (.Y (nx10396), .A0 (nx29069), .A1 (nx34419), .B0 (nx29073)) ;
    dffr reg_label_5_input_state_machine_0 (.Q (label_5_input_state_machine_0), 
         .QB (nx29069), .D (nx20183), .CLK (clk), .R (rst)) ;
    oai21 ix29074 (.Y (nx29073), .A0 (nx35763), .A1 (label_5_output[0]), .B0 (
          nx10384)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_4_1), .QB (\$dummy [286]), .D (nx20163)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_4_2), .QB (nx29494), .D (nx20153), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_4_3), .QB (\$dummy [287]), .D (nx20143)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_4_4), .QB (nx29492), .D (nx20133), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_4_5), .QB (\$dummy [288]), .D (nx20123)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_4_6), .QB (nx29490), .D (nx20113), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_4_7), .QB (\$dummy [289]), .D (nx20103)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_4_8), .QB (nx29488), .D (nx20093), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_4_9), .QB (\$dummy [290]), .D (nx20083)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_4_10), .QB (nx29486), .D (nx20073), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_4_11), .QB (\$dummy [291]), .D (nx20063)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_4_12), .QB (nx29484), .D (nx20053), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_4_13), .QB (\$dummy [292]), .D (nx20043)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_4_14), .QB (nx29482), .D (nx20033), .CLK (
         clk), .R (rst)) ;
    aoi22 ix29123 (.Y (nx29122), .A0 (mdr_data_out[15]), .A1 (nx34939), .B0 (
          nx10182), .B1 (nx10188)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_reg_output_0), .QB (\$dummy [293]), .D (
         nx19673), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_4_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_4_shift_Reg_count_0), .QB (\$dummy [294]), .D (
            nx19659), .CLK (clk), .S (nx34481)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_reg_output_9), .QB (\$dummy [295]), .D (
         nx19853), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_9), .QB (\$dummy [296]), .D (
         nx19843), .CLK (clk), .R (nx34481)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_8), .QB (\$dummy [297]), .D (
         nx19833), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_8), .QB (\$dummy [298]), .D (
         nx19823), .CLK (clk), .R (nx34479)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_7), .QB (\$dummy [299]), .D (
         nx19813), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_7), .QB (\$dummy [300]), .D (
         nx19803), .CLK (clk), .R (nx34479)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_6), .QB (\$dummy [301]), .D (
         nx19793), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_6), .QB (\$dummy [302]), .D (
         nx19783), .CLK (clk), .R (nx34479)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_5), .QB (\$dummy [303]), .D (
         nx19773), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_5), .QB (\$dummy [304]), .D (
         nx19763), .CLK (clk), .R (nx34479)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_4), .QB (\$dummy [305]), .D (
         nx19753), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_4), .QB (\$dummy [306]), .D (
         nx19743), .CLK (clk), .R (nx34479)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_3), .QB (\$dummy [307]), .D (
         nx19733), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_3), .QB (\$dummy [308]), .D (
         nx19723), .CLK (clk), .R (nx34479)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_2), .QB (\$dummy [309]), .D (
         nx19713), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_2), .QB (\$dummy [310]), .D (
         nx19703), .CLK (clk), .R (nx34479)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_4_shift_Reg_output_1), .QB (\$dummy [311]), .D (
         nx19693), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_4_shift_Reg_count_1), .QB (\$dummy [312]), .D (
         nx19683), .CLK (clk), .R (nx34477)) ;
    nand02 ix19654 (.Y (nx19653), .A0 (nx35823), .A1 (nx34925)) ;
    dffs_ni booth_booth_integrtaion_4_shift_Reg_reg_en (.Q (\$dummy [313]), .QB (
            nx29169), .D (nx19653), .CLK (clk), .S (nx34477)) ;
    nand02 ix10183 (.Y (nx10182), .A0 (nx29190), .A1 (nx29202)) ;
    oai21 ix29191 (.Y (nx29190), .A0 (nx34953), .A1 (nx34947), .B0 (
          mdr_data_out[80])) ;
    oai21 ix19864 (.Y (nx19863), .A0 (nx29195), .A1 (nx35425), .B0 (nx29197)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [314]), .QB (
         nx29195), .D (nx19863), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [315]), .QB (
         nx29199), .D (nx20173), .CLK (clk), .R (rst)) ;
    xnor2 ix29207 (.Y (nx29206), .A0 (nx9652), .A1 (nx13217)) ;
    oai21 ix20004 (.Y (nx20003), .A0 (nx29212), .A1 (nx35425), .B0 (nx29214)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_17), .QB (nx29212), .D (nx20003)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29215 (.Y (nx29214), .A0 (nx35433), .A1 (nx10160), .A2 (nx36109)) ;
    xnor2 ix10161 (.Y (nx10160), .A0 (nx29217), .A1 (nx13219)) ;
    aoi22 ix29218 (.Y (nx29217), .A0 (booth_booth_integrtaion_4_booth_output_17)
          , .A1 (nx9676), .B0 (nx9652), .B1 (nx13217)) ;
    nand02 ix9661 (.Y (nx9660), .A0 (mdr_data_out[81]), .A1 (mdr_data_out[80])
           ) ;
    or02 ix29222 (.Y (nx29221), .A0 (mdr_data_out[80]), .A1 (mdr_data_out[81])
         ) ;
    xnor2 ix29228 (.Y (nx29227), .A0 (nx9704), .A1 (nx13221)) ;
    oai22 ix9705 (.Y (nx9704), .A0 (nx29217), .A1 (nx29230), .B0 (nx29237), .B1 (
          nx35437)) ;
    aoi32 ix29233 (.Y (nx29232), .A0 (nx9686), .A1 (nx34953), .A2 (nx29235), .B0 (
          mdr_data_out[82]), .B1 (nx34947)) ;
    oai21 ix9687 (.Y (nx9686), .A0 (mdr_data_out[80]), .A1 (mdr_data_out[81]), .B0 (
          mdr_data_out[82])) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_18), .QB (nx29237), .D (nx19993)
         , .CLK (clk), .R (rst)) ;
    oai21 ix19984 (.Y (nx19983), .A0 (nx29242), .A1 (nx35425), .B0 (nx29244)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_19), .QB (nx29242), .D (nx19983)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29245 (.Y (nx29244), .A0 (nx35433), .A1 (nx10136), .A2 (nx36109)) ;
    xnor2 ix10137 (.Y (nx10136), .A0 (nx29247), .A1 (nx13223)) ;
    aoi22 ix29248 (.Y (nx29247), .A0 (booth_booth_integrtaion_4_booth_output_19)
          , .A1 (nx9724), .B0 (nx9704), .B1 (nx13221)) ;
    nor02ii ix29251 (.Y (nx29250), .A0 (nx9690), .A1 (mdr_data_out[83])) ;
    nor03_2x ix9691 (.Y (nx9690), .A0 (mdr_data_out[82]), .A1 (mdr_data_out[80])
             , .A2 (mdr_data_out[81])) ;
    nor04 ix9715 (.Y (nx9714), .A0 (mdr_data_out[83]), .A1 (mdr_data_out[82]), .A2 (
          mdr_data_out[80]), .A3 (mdr_data_out[81])) ;
    xnor2 ix29265 (.Y (nx29264), .A0 (nx9752), .A1 (nx13224)) ;
    oai22 ix9753 (.Y (nx9752), .A0 (nx29247), .A1 (nx29267), .B0 (nx29276), .B1 (
          nx35439)) ;
    aoi32 ix29270 (.Y (nx29269), .A0 (nx9734), .A1 (nx34953), .A2 (nx29274), .B0 (
          mdr_data_out[84]), .B1 (nx34947)) ;
    nand02 ix9735 (.Y (nx9734), .A0 (nx29272), .A1 (mdr_data_out[84])) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_20), .QB (nx29276), .D (nx19973)
         , .CLK (clk), .R (rst)) ;
    oai21 ix19964 (.Y (nx19963), .A0 (nx29281), .A1 (nx35425), .B0 (nx29283)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_21), .QB (nx29281), .D (nx19963)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29284 (.Y (nx29283), .A0 (nx35433), .A1 (nx10112), .A2 (nx36109)) ;
    xnor2 ix10113 (.Y (nx10112), .A0 (nx29286), .A1 (nx13225)) ;
    aoi22 ix29287 (.Y (nx29286), .A0 (booth_booth_integrtaion_4_booth_output_21)
          , .A1 (nx9772), .B0 (nx9752), .B1 (nx13224)) ;
    nor02ii ix29290 (.Y (nx29289), .A0 (nx9738), .A1 (mdr_data_out[85])) ;
    nor02ii ix9739 (.Y (nx9738), .A0 (mdr_data_out[84]), .A1 (nx9714)) ;
    nor02ii ix9763 (.Y (nx9762), .A0 (mdr_data_out[85]), .A1 (nx9738)) ;
    xnor2 ix29300 (.Y (nx29299), .A0 (nx9800), .A1 (nx13226)) ;
    oai22 ix9801 (.Y (nx9800), .A0 (nx29286), .A1 (nx29302), .B0 (nx29311), .B1 (
          nx35441)) ;
    aoi32 ix29305 (.Y (nx29304), .A0 (nx9782), .A1 (nx34953), .A2 (nx29309), .B0 (
          mdr_data_out[86]), .B1 (nx34947)) ;
    nand02 ix9783 (.Y (nx9782), .A0 (nx29307), .A1 (mdr_data_out[86])) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_22), .QB (nx29311), .D (nx19953)
         , .CLK (clk), .R (rst)) ;
    oai21 ix19944 (.Y (nx19943), .A0 (nx29316), .A1 (nx35425), .B0 (nx29318)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_23), .QB (nx29316), .D (nx19943)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29319 (.Y (nx29318), .A0 (nx35433), .A1 (nx10088), .A2 (nx35427)) ;
    xnor2 ix10089 (.Y (nx10088), .A0 (nx29321), .A1 (nx13227)) ;
    aoi22 ix29322 (.Y (nx29321), .A0 (booth_booth_integrtaion_4_booth_output_23)
          , .A1 (nx9820), .B0 (nx9800), .B1 (nx13226)) ;
    nor02ii ix29325 (.Y (nx29324), .A0 (nx9786), .A1 (mdr_data_out[87])) ;
    nor02ii ix9787 (.Y (nx9786), .A0 (mdr_data_out[86]), .A1 (nx9762)) ;
    nor02ii ix9811 (.Y (nx9810), .A0 (mdr_data_out[87]), .A1 (nx9786)) ;
    xnor2 ix29335 (.Y (nx29334), .A0 (nx9848), .A1 (nx13228)) ;
    oai22 ix9849 (.Y (nx9848), .A0 (nx29321), .A1 (nx29337), .B0 (nx29346), .B1 (
          nx35443)) ;
    aoi32 ix29340 (.Y (nx29339), .A0 (nx9830), .A1 (nx34953), .A2 (nx29344), .B0 (
          mdr_data_out[88]), .B1 (nx34947)) ;
    nand02 ix9831 (.Y (nx9830), .A0 (nx29342), .A1 (mdr_data_out[88])) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_24), .QB (nx29346), .D (nx19933)
         , .CLK (clk), .R (rst)) ;
    oai21 ix19924 (.Y (nx19923), .A0 (nx29351), .A1 (nx35427), .B0 (nx29353)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_25), .QB (nx29351), .D (nx19923)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29354 (.Y (nx29353), .A0 (nx35433), .A1 (nx10064), .A2 (nx35427)) ;
    xnor2 ix10065 (.Y (nx10064), .A0 (nx29356), .A1 (nx13229)) ;
    aoi22 ix29357 (.Y (nx29356), .A0 (booth_booth_integrtaion_4_booth_output_25)
          , .A1 (nx9868), .B0 (nx9848), .B1 (nx13228)) ;
    nor02ii ix29360 (.Y (nx29359), .A0 (nx9834), .A1 (mdr_data_out[89])) ;
    nor02ii ix9835 (.Y (nx9834), .A0 (mdr_data_out[88]), .A1 (nx9810)) ;
    nor02ii ix9859 (.Y (nx9858), .A0 (mdr_data_out[89]), .A1 (nx9834)) ;
    xnor2 ix29370 (.Y (nx29369), .A0 (nx9896), .A1 (nx13231)) ;
    oai22 ix9897 (.Y (nx9896), .A0 (nx29356), .A1 (nx29372), .B0 (nx29381), .B1 (
          nx35445)) ;
    aoi32 ix29375 (.Y (nx29374), .A0 (nx9878), .A1 (nx34953), .A2 (nx29379), .B0 (
          mdr_data_out[90]), .B1 (nx34947)) ;
    nand02 ix9879 (.Y (nx9878), .A0 (nx29377), .A1 (mdr_data_out[90])) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_26), .QB (nx29381), .D (nx19913)
         , .CLK (clk), .R (rst)) ;
    oai21 ix19904 (.Y (nx19903), .A0 (nx29386), .A1 (nx35427), .B0 (nx29388)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_27), .QB (nx29386), .D (nx19903)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29389 (.Y (nx29388), .A0 (nx35433), .A1 (nx10040), .A2 (nx35427)) ;
    xnor2 ix10041 (.Y (nx10040), .A0 (nx29391), .A1 (nx13233)) ;
    aoi22 ix29392 (.Y (nx29391), .A0 (booth_booth_integrtaion_4_booth_output_27)
          , .A1 (nx9916), .B0 (nx9896), .B1 (nx13231)) ;
    nor02ii ix29395 (.Y (nx29394), .A0 (nx9882), .A1 (mdr_data_out[91])) ;
    nor02ii ix9883 (.Y (nx9882), .A0 (mdr_data_out[90]), .A1 (nx9858)) ;
    nor02ii ix9907 (.Y (nx9906), .A0 (mdr_data_out[91]), .A1 (nx9882)) ;
    xnor2 ix29405 (.Y (nx29404), .A0 (nx9944), .A1 (nx13235)) ;
    oai22 ix9945 (.Y (nx9944), .A0 (nx29391), .A1 (nx29407), .B0 (nx29416), .B1 (
          nx35447)) ;
    aoi32 ix29410 (.Y (nx29409), .A0 (nx9926), .A1 (nx34953), .A2 (nx29414), .B0 (
          mdr_data_out[92]), .B1 (nx34947)) ;
    nand02 ix9927 (.Y (nx9926), .A0 (nx29412), .A1 (mdr_data_out[92])) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_28), .QB (nx29416), .D (nx19893)
         , .CLK (clk), .R (rst)) ;
    oai21 ix19884 (.Y (nx19883), .A0 (nx29421), .A1 (nx35427), .B0 (nx29423)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_29), .QB (nx29421), .D (nx19883)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29424 (.Y (nx29423), .A0 (nx36117), .A1 (nx10016), .A2 (nx35427)) ;
    xnor2 ix10017 (.Y (nx10016), .A0 (nx29426), .A1 (nx13236)) ;
    aoi22 ix29427 (.Y (nx29426), .A0 (booth_booth_integrtaion_4_booth_output_29)
          , .A1 (nx9964), .B0 (nx9944), .B1 (nx13235)) ;
    nor02ii ix29430 (.Y (nx29429), .A0 (nx9930), .A1 (mdr_data_out[93])) ;
    nor02ii ix9931 (.Y (nx9930), .A0 (mdr_data_out[92]), .A1 (nx9906)) ;
    nor02ii ix9955 (.Y (nx9954), .A0 (mdr_data_out[93]), .A1 (nx9930)) ;
    xnor2 ix29440 (.Y (nx29439), .A0 (nx9992), .A1 (nx10002)) ;
    oai22 ix9993 (.Y (nx9992), .A0 (nx29426), .A1 (nx29442), .B0 (nx29451), .B1 (
          nx35449)) ;
    aoi32 ix29445 (.Y (nx29444), .A0 (nx9974), .A1 (nx34955), .A2 (nx29449), .B0 (
          mdr_data_out[94]), .B1 (nx34949)) ;
    nand02 ix9975 (.Y (nx9974), .A0 (nx29447), .A1 (mdr_data_out[94])) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_31), .QB (nx29451), .D (nx19873)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix29455 (.Y (nx29454), .A0 (mdr_data_out[95]), .A1 (nx34949), .B0 (
          nx34955), .B1 (nx9994)) ;
    xnor2 ix9995 (.Y (nx9994), .A0 (mdr_data_out[95]), .A1 (nx9978)) ;
    nor02ii ix9979 (.Y (nx9978), .A0 (mdr_data_out[94]), .A1 (nx9954)) ;
    aoi32 ix29459 (.Y (nx29458), .A0 (nx9950), .A1 (nx34955), .A2 (nx29447), .B0 (
          mdr_data_out[93]), .B1 (nx34949)) ;
    aoi32 ix29462 (.Y (nx29461), .A0 (nx9902), .A1 (nx34955), .A2 (nx29412), .B0 (
          mdr_data_out[91]), .B1 (nx34949)) ;
    aoi32 ix29465 (.Y (nx29464), .A0 (nx9854), .A1 (nx34955), .A2 (nx29377), .B0 (
          mdr_data_out[89]), .B1 (nx34949)) ;
    aoi32 ix29468 (.Y (nx29467), .A0 (nx9806), .A1 (nx34955), .A2 (nx29342), .B0 (
          mdr_data_out[87]), .B1 (nx34949)) ;
    aoi32 ix29471 (.Y (nx29470), .A0 (nx9758), .A1 (nx34955), .A2 (nx29307), .B0 (
          mdr_data_out[85]), .B1 (nx34949)) ;
    aoi32 ix29474 (.Y (nx29473), .A0 (nx9710), .A1 (nx9646), .A2 (nx29272), .B0 (
          mdr_data_out[83]), .B1 (nx34951)) ;
    aoi32 ix29477 (.Y (nx29476), .A0 (nx9660), .A1 (nx9646), .A2 (nx29221), .B0 (
          mdr_data_out[81]), .B1 (nx34951)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_4_booth_output_16), .QB (nx29202), .D (nx20013)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_4_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_4_15), .QB (nx29480), .D (nx20023), .CLK (
         clk), .R (rst)) ;
    aoi21 ix10385 (.Y (nx10384), .A0 (label_5_output[0]), .A1 (nx35763), .B0 (
          nx36387)) ;
    oai21 ix21584 (.Y (nx21583), .A0 (nx29502), .A1 (nx34765), .B0 (nx29504)) ;
    dff max_calc_reg_comparator_third_inp2_0 (.Q (\$dummy [316]), .QB (nx29502)
        , .D (nx21583), .CLK (clk)) ;
    nand03 ix29505 (.Y (nx29504), .A0 (label_6_output[0]), .A1 (nx35453), .A2 (
           nx34765)) ;
    dffr labelsregfile_label6_loop1_0_fx_reg_q (.Q (label_6_output[0]), .QB (
         \$dummy [317]), .D (nx21033), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_0 (.Q (label_6_input_0), .D (nx11718), .CLK (nx34521
          )) ;
    oai21 ix11719 (.Y (nx11718), .A0 (nx29510), .A1 (nx34419), .B0 (nx29514)) ;
    dffr reg_label_6_input_state_machine_0 (.Q (label_6_input_state_machine_0), 
         .QB (nx29510), .D (nx21023), .CLK (clk), .R (rst)) ;
    oai21 ix29515 (.Y (nx29514), .A0 (nx35767), .A1 (label_6_output[0]), .B0 (
          nx11706)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_5_1), .QB (\$dummy [318]), .D (nx21003)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_5_2), .QB (nx29935), .D (nx20993), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_5_3), .QB (\$dummy [319]), .D (nx20983)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_5_4), .QB (nx29933), .D (nx20973), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_5_5), .QB (\$dummy [320]), .D (nx20963)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_5_6), .QB (nx29931), .D (nx20953), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_5_7), .QB (\$dummy [321]), .D (nx20943)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_5_8), .QB (nx29929), .D (nx20933), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_5_9), .QB (\$dummy [322]), .D (nx20923)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_5_10), .QB (nx29927), .D (nx20913), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_5_11), .QB (\$dummy [323]), .D (nx20903)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_5_12), .QB (nx29925), .D (nx20893), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_5_13), .QB (\$dummy [324]), .D (nx20883)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_5_14), .QB (nx29923), .D (nx20873), .CLK (
         clk), .R (rst)) ;
    aoi22 ix29564 (.Y (nx29563), .A0 (mdr_data_out[15]), .A1 (nx34971), .B0 (
          nx11504), .B1 (nx11510)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_reg_output_0), .QB (\$dummy [325]), .D (
         nx20513), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_5_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_5_shift_Reg_count_0), .QB (\$dummy [326]), .D (
            nx20499), .CLK (clk), .S (nx34483)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_reg_output_9), .QB (\$dummy [327]), .D (
         nx20693), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_9), .QB (\$dummy [328]), .D (
         nx20683), .CLK (clk), .R (nx34483)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_8), .QB (\$dummy [329]), .D (
         nx20673), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_8), .QB (\$dummy [330]), .D (
         nx20663), .CLK (clk), .R (nx34483)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_7), .QB (\$dummy [331]), .D (
         nx20653), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_7), .QB (\$dummy [332]), .D (
         nx20643), .CLK (clk), .R (nx34483)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_6), .QB (\$dummy [333]), .D (
         nx20633), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_6), .QB (\$dummy [334]), .D (
         nx20623), .CLK (clk), .R (nx34483)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_5), .QB (\$dummy [335]), .D (
         nx20613), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_5), .QB (\$dummy [336]), .D (
         nx20603), .CLK (clk), .R (nx34483)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_4), .QB (\$dummy [337]), .D (
         nx20593), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_4), .QB (\$dummy [338]), .D (
         nx20583), .CLK (clk), .R (nx34481)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_3), .QB (\$dummy [339]), .D (
         nx20573), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_3), .QB (\$dummy [340]), .D (
         nx20563), .CLK (clk), .R (nx34481)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_2), .QB (\$dummy [341]), .D (
         nx20553), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_2), .QB (\$dummy [342]), .D (
         nx20543), .CLK (clk), .R (nx34481)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_5_shift_Reg_output_1), .QB (\$dummy [343]), .D (
         nx20533), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_5_shift_Reg_count_1), .QB (\$dummy [344]), .D (
         nx20523), .CLK (clk), .R (nx34481)) ;
    nand02 ix20494 (.Y (nx20493), .A0 (nx35827), .A1 (nx34957)) ;
    dffs_ni booth_booth_integrtaion_5_shift_Reg_reg_en (.Q (\$dummy [345]), .QB (
            nx29610), .D (nx20493), .CLK (clk), .S (nx34481)) ;
    nand02 ix11505 (.Y (nx11504), .A0 (nx29631), .A1 (nx29643)) ;
    oai21 ix29632 (.Y (nx29631), .A0 (nx34985), .A1 (nx34979), .B0 (
          mdr_data_out[96])) ;
    oai21 ix20704 (.Y (nx20703), .A0 (nx29636), .A1 (nx35473), .B0 (nx29638)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [346]), .QB (
         nx29636), .D (nx20703), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [347]), .QB (
         nx29640), .D (nx21013), .CLK (clk), .R (rst)) ;
    xnor2 ix29648 (.Y (nx29647), .A0 (nx10974), .A1 (nx13257)) ;
    oai21 ix20844 (.Y (nx20843), .A0 (nx29653), .A1 (nx35473), .B0 (nx29655)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_17), .QB (nx29653), .D (nx20843)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29656 (.Y (nx29655), .A0 (nx35481), .A1 (nx11482), .A2 (nx36131)) ;
    xnor2 ix11483 (.Y (nx11482), .A0 (nx29658), .A1 (nx13259)) ;
    aoi22 ix29659 (.Y (nx29658), .A0 (booth_booth_integrtaion_5_booth_output_17)
          , .A1 (nx10998), .B0 (nx10974), .B1 (nx13257)) ;
    nand02 ix10983 (.Y (nx10982), .A0 (mdr_data_out[97]), .A1 (mdr_data_out[96])
           ) ;
    or02 ix29663 (.Y (nx29662), .A0 (mdr_data_out[96]), .A1 (mdr_data_out[97])
         ) ;
    xnor2 ix29669 (.Y (nx29668), .A0 (nx11026), .A1 (nx13260)) ;
    oai22 ix11027 (.Y (nx11026), .A0 (nx29658), .A1 (nx29671), .B0 (nx29678), .B1 (
          nx35485)) ;
    aoi32 ix29674 (.Y (nx29673), .A0 (nx11008), .A1 (nx34985), .A2 (nx29676), .B0 (
          mdr_data_out[98]), .B1 (nx34979)) ;
    oai21 ix11009 (.Y (nx11008), .A0 (mdr_data_out[96]), .A1 (mdr_data_out[97])
          , .B0 (mdr_data_out[98])) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_18), .QB (nx29678), .D (nx20833)
         , .CLK (clk), .R (rst)) ;
    oai21 ix20824 (.Y (nx20823), .A0 (nx29683), .A1 (nx35473), .B0 (nx29685)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_19), .QB (nx29683), .D (nx20823)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29686 (.Y (nx29685), .A0 (nx35481), .A1 (nx11458), .A2 (nx36131)) ;
    xnor2 ix11459 (.Y (nx11458), .A0 (nx29688), .A1 (nx13261)) ;
    aoi22 ix29689 (.Y (nx29688), .A0 (booth_booth_integrtaion_5_booth_output_19)
          , .A1 (nx11046), .B0 (nx11026), .B1 (nx13260)) ;
    nor02ii ix29692 (.Y (nx29691), .A0 (nx11012), .A1 (mdr_data_out[99])) ;
    nor03_2x ix11013 (.Y (nx11012), .A0 (mdr_data_out[98]), .A1 (
             mdr_data_out[96]), .A2 (mdr_data_out[97])) ;
    nor04 ix11037 (.Y (nx11036), .A0 (mdr_data_out[99]), .A1 (mdr_data_out[98])
          , .A2 (mdr_data_out[96]), .A3 (mdr_data_out[97])) ;
    xnor2 ix29706 (.Y (nx29705), .A0 (nx11074), .A1 (nx13262)) ;
    oai22 ix11075 (.Y (nx11074), .A0 (nx29688), .A1 (nx29708), .B0 (nx29717), .B1 (
          nx35487)) ;
    aoi32 ix29711 (.Y (nx29710), .A0 (nx11056), .A1 (nx34985), .A2 (nx29715), .B0 (
          mdr_data_out[100]), .B1 (nx34979)) ;
    nand02 ix11057 (.Y (nx11056), .A0 (nx29713), .A1 (mdr_data_out[100])) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_20), .QB (nx29717), .D (nx20813)
         , .CLK (clk), .R (rst)) ;
    oai21 ix20804 (.Y (nx20803), .A0 (nx29722), .A1 (nx35473), .B0 (nx29724)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_21), .QB (nx29722), .D (nx20803)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29725 (.Y (nx29724), .A0 (nx35481), .A1 (nx11434), .A2 (nx36131)) ;
    xnor2 ix11435 (.Y (nx11434), .A0 (nx29727), .A1 (nx13263)) ;
    aoi22 ix29728 (.Y (nx29727), .A0 (booth_booth_integrtaion_5_booth_output_21)
          , .A1 (nx11094), .B0 (nx11074), .B1 (nx13262)) ;
    nor02ii ix29731 (.Y (nx29730), .A0 (nx11060), .A1 (mdr_data_out[101])) ;
    nor02ii ix11061 (.Y (nx11060), .A0 (mdr_data_out[100]), .A1 (nx11036)) ;
    nor02ii ix11085 (.Y (nx11084), .A0 (mdr_data_out[101]), .A1 (nx11060)) ;
    xnor2 ix29741 (.Y (nx29740), .A0 (nx11122), .A1 (nx13264)) ;
    oai22 ix11123 (.Y (nx11122), .A0 (nx29727), .A1 (nx29743), .B0 (nx29752), .B1 (
          nx35489)) ;
    aoi32 ix29746 (.Y (nx29745), .A0 (nx11104), .A1 (nx34985), .A2 (nx29750), .B0 (
          mdr_data_out[102]), .B1 (nx34979)) ;
    nand02 ix11105 (.Y (nx11104), .A0 (nx29748), .A1 (mdr_data_out[102])) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_22), .QB (nx29752), .D (nx20793)
         , .CLK (clk), .R (rst)) ;
    oai21 ix20784 (.Y (nx20783), .A0 (nx29757), .A1 (nx35473), .B0 (nx29759)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_23), .QB (nx29757), .D (nx20783)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29760 (.Y (nx29759), .A0 (nx35481), .A1 (nx11410), .A2 (nx35475)) ;
    xnor2 ix11411 (.Y (nx11410), .A0 (nx29762), .A1 (nx13265)) ;
    aoi22 ix29763 (.Y (nx29762), .A0 (booth_booth_integrtaion_5_booth_output_23)
          , .A1 (nx11142), .B0 (nx11122), .B1 (nx13264)) ;
    nor02ii ix29766 (.Y (nx29765), .A0 (nx11108), .A1 (mdr_data_out[103])) ;
    nor02ii ix11109 (.Y (nx11108), .A0 (mdr_data_out[102]), .A1 (nx11084)) ;
    nor02ii ix11133 (.Y (nx11132), .A0 (mdr_data_out[103]), .A1 (nx11108)) ;
    xnor2 ix29776 (.Y (nx29775), .A0 (nx11170), .A1 (nx13267)) ;
    oai22 ix11171 (.Y (nx11170), .A0 (nx29762), .A1 (nx29778), .B0 (nx29787), .B1 (
          nx35491)) ;
    aoi32 ix29781 (.Y (nx29780), .A0 (nx11152), .A1 (nx34985), .A2 (nx29785), .B0 (
          mdr_data_out[104]), .B1 (nx34979)) ;
    nand02 ix11153 (.Y (nx11152), .A0 (nx29783), .A1 (mdr_data_out[104])) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_24), .QB (nx29787), .D (nx20773)
         , .CLK (clk), .R (rst)) ;
    oai21 ix20764 (.Y (nx20763), .A0 (nx29792), .A1 (nx35475), .B0 (nx29794)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_25), .QB (nx29792), .D (nx20763)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29795 (.Y (nx29794), .A0 (nx35481), .A1 (nx11386), .A2 (nx35475)) ;
    xnor2 ix11387 (.Y (nx11386), .A0 (nx29797), .A1 (nx13269)) ;
    aoi22 ix29798 (.Y (nx29797), .A0 (booth_booth_integrtaion_5_booth_output_25)
          , .A1 (nx11190), .B0 (nx11170), .B1 (nx13267)) ;
    nor02ii ix29801 (.Y (nx29800), .A0 (nx11156), .A1 (mdr_data_out[105])) ;
    nor02ii ix11157 (.Y (nx11156), .A0 (mdr_data_out[104]), .A1 (nx11132)) ;
    nor02ii ix11181 (.Y (nx11180), .A0 (mdr_data_out[105]), .A1 (nx11156)) ;
    xnor2 ix29811 (.Y (nx29810), .A0 (nx11218), .A1 (nx13271)) ;
    oai22 ix11219 (.Y (nx11218), .A0 (nx29797), .A1 (nx29813), .B0 (nx29822), .B1 (
          nx35493)) ;
    aoi32 ix29816 (.Y (nx29815), .A0 (nx11200), .A1 (nx34985), .A2 (nx29820), .B0 (
          mdr_data_out[106]), .B1 (nx34979)) ;
    nand02 ix11201 (.Y (nx11200), .A0 (nx29818), .A1 (mdr_data_out[106])) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_26), .QB (nx29822), .D (nx20753)
         , .CLK (clk), .R (rst)) ;
    oai21 ix20744 (.Y (nx20743), .A0 (nx29827), .A1 (nx35475), .B0 (nx29829)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_27), .QB (nx29827), .D (nx20743)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29830 (.Y (nx29829), .A0 (nx35481), .A1 (nx11362), .A2 (nx35475)) ;
    xnor2 ix11363 (.Y (nx11362), .A0 (nx29832), .A1 (nx13272)) ;
    aoi22 ix29833 (.Y (nx29832), .A0 (booth_booth_integrtaion_5_booth_output_27)
          , .A1 (nx11238), .B0 (nx11218), .B1 (nx13271)) ;
    nor02ii ix29836 (.Y (nx29835), .A0 (nx11204), .A1 (mdr_data_out[107])) ;
    nor02ii ix11205 (.Y (nx11204), .A0 (mdr_data_out[106]), .A1 (nx11180)) ;
    nor02ii ix11229 (.Y (nx11228), .A0 (mdr_data_out[107]), .A1 (nx11204)) ;
    xnor2 ix29846 (.Y (nx29845), .A0 (nx11266), .A1 (nx13273)) ;
    oai22 ix11267 (.Y (nx11266), .A0 (nx29832), .A1 (nx29848), .B0 (nx29857), .B1 (
          nx35495)) ;
    aoi32 ix29851 (.Y (nx29850), .A0 (nx11248), .A1 (nx34985), .A2 (nx29855), .B0 (
          mdr_data_out[108]), .B1 (nx34979)) ;
    nand02 ix11249 (.Y (nx11248), .A0 (nx29853), .A1 (mdr_data_out[108])) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_28), .QB (nx29857), .D (nx20733)
         , .CLK (clk), .R (rst)) ;
    oai21 ix20724 (.Y (nx20723), .A0 (nx29862), .A1 (nx35475), .B0 (nx29864)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_29), .QB (nx29862), .D (nx20723)
         , .CLK (clk), .R (rst)) ;
    nand03 ix29865 (.Y (nx29864), .A0 (nx36139), .A1 (nx11338), .A2 (nx35475)) ;
    xnor2 ix11339 (.Y (nx11338), .A0 (nx29867), .A1 (nx13274)) ;
    aoi22 ix29868 (.Y (nx29867), .A0 (booth_booth_integrtaion_5_booth_output_29)
          , .A1 (nx11286), .B0 (nx11266), .B1 (nx13273)) ;
    nor02ii ix29871 (.Y (nx29870), .A0 (nx11252), .A1 (mdr_data_out[109])) ;
    nor02ii ix11253 (.Y (nx11252), .A0 (mdr_data_out[108]), .A1 (nx11228)) ;
    nor02ii ix11277 (.Y (nx11276), .A0 (mdr_data_out[109]), .A1 (nx11252)) ;
    xnor2 ix29881 (.Y (nx29880), .A0 (nx11314), .A1 (nx11324)) ;
    oai22 ix11315 (.Y (nx11314), .A0 (nx29867), .A1 (nx29883), .B0 (nx29892), .B1 (
          nx35497)) ;
    aoi32 ix29886 (.Y (nx29885), .A0 (nx11296), .A1 (nx34987), .A2 (nx29890), .B0 (
          mdr_data_out[110]), .B1 (nx34981)) ;
    nand02 ix11297 (.Y (nx11296), .A0 (nx29888), .A1 (mdr_data_out[110])) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_31), .QB (nx29892), .D (nx20713)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix29896 (.Y (nx29895), .A0 (mdr_data_out[111]), .A1 (nx34981), .B0 (
          nx34987), .B1 (nx11316)) ;
    xnor2 ix11317 (.Y (nx11316), .A0 (mdr_data_out[111]), .A1 (nx11300)) ;
    nor02ii ix11301 (.Y (nx11300), .A0 (mdr_data_out[110]), .A1 (nx11276)) ;
    aoi32 ix29900 (.Y (nx29899), .A0 (nx11272), .A1 (nx34987), .A2 (nx29888), .B0 (
          mdr_data_out[109]), .B1 (nx34981)) ;
    aoi32 ix29903 (.Y (nx29902), .A0 (nx11224), .A1 (nx34987), .A2 (nx29853), .B0 (
          mdr_data_out[107]), .B1 (nx34981)) ;
    aoi32 ix29906 (.Y (nx29905), .A0 (nx11176), .A1 (nx34987), .A2 (nx29818), .B0 (
          mdr_data_out[105]), .B1 (nx34981)) ;
    aoi32 ix29909 (.Y (nx29908), .A0 (nx11128), .A1 (nx34987), .A2 (nx29783), .B0 (
          mdr_data_out[103]), .B1 (nx34981)) ;
    aoi32 ix29912 (.Y (nx29911), .A0 (nx11080), .A1 (nx34987), .A2 (nx29748), .B0 (
          mdr_data_out[101]), .B1 (nx34981)) ;
    aoi32 ix29915 (.Y (nx29914), .A0 (nx11032), .A1 (nx10968), .A2 (nx29713), .B0 (
          mdr_data_out[99]), .B1 (nx34983)) ;
    aoi32 ix29918 (.Y (nx29917), .A0 (nx10982), .A1 (nx10968), .A2 (nx29662), .B0 (
          mdr_data_out[97]), .B1 (nx34983)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_5_booth_output_16), .QB (nx29643), .D (nx20853)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_5_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_5_15), .QB (nx29921), .D (nx20863), .CLK (
         clk), .R (rst)) ;
    aoi21 ix11707 (.Y (nx11706), .A0 (label_6_output[0]), .A1 (nx35767), .B0 (
          nx36387)) ;
    xnor2 ix12691 (.Y (nx12690), .A0 (nx29940), .A1 (nx12688)) ;
    aoi22 ix29941 (.Y (nx29940), .A0 (nx29942), .A1 (
          max_calc_comparator_third_inp1_14), .B0 (nx12176), .B1 (nx12594)) ;
    dff max_calc_reg_comparator_third_inp2_14 (.Q (\$dummy [348]), .QB (nx29942)
        , .D (nx21313), .CLK (clk)) ;
    oai21 ix21314 (.Y (nx21313), .A0 (nx29942), .A1 (nx34765), .B0 (nx29945)) ;
    dffr labelsregfile_label6_loop1_14_fx_reg_q (.Q (label_6_output[14]), .QB (
         nx30129), .D (nx21303), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_14 (.Q (label_6_input_14), .D (nx12154), .CLK (
          nx34525)) ;
    dffr reg_label_6_input_state_machine_14 (.Q (label_6_input_state_machine_14)
         , .QB (\$dummy [349]), .D (nx20483), .CLK (clk), .R (rst)) ;
    xor2 ix12151 (.Y (nx12150), .A0 (nx29955), .A1 (nx30127)) ;
    aoi22 ix29956 (.Y (nx29955), .A0 (label_6_output[13]), .A1 (
          booth_booth_integration_output_5_13), .B0 (nx12114), .B1 (nx13293)) ;
    dffr labelsregfile_label6_loop1_13_fx_reg_q (.Q (label_6_output[13]), .QB (
         \$dummy [350]), .D (nx21293), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_13 (.Q (label_6_input_13), .D (nx12128), .CLK (
          nx34525)) ;
    dffr reg_label_6_input_state_machine_13 (.Q (label_6_input_state_machine_13)
         , .QB (\$dummy [351]), .D (nx21283), .CLK (clk), .R (rst)) ;
    xnor2 ix12125 (.Y (nx12124), .A0 (nx12114), .A1 (nx30123)) ;
    oai22 ix12115 (.Y (nx12114), .A0 (nx29966), .A1 (nx30112), .B0 (nx30122), .B1 (
          nx29925)) ;
    aoi22 ix29967 (.Y (nx29966), .A0 (label_6_output[11]), .A1 (
          booth_booth_integration_output_5_11), .B0 (nx12050), .B1 (nx13289)) ;
    dffr labelsregfile_label6_loop1_11_fx_reg_q (.Q (label_6_output[11]), .QB (
         \$dummy [352]), .D (nx21253), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_11 (.Q (label_6_input_11), .D (nx12064), .CLK (
          nx34523)) ;
    dffr reg_label_6_input_state_machine_11 (.Q (label_6_input_state_machine_11)
         , .QB (\$dummy [353]), .D (nx21243), .CLK (clk), .R (rst)) ;
    xnor2 ix12061 (.Y (nx12060), .A0 (nx12050), .A1 (nx30108)) ;
    oai22 ix12051 (.Y (nx12050), .A0 (nx29977), .A1 (nx30097), .B0 (nx30107), .B1 (
          nx29927)) ;
    aoi22 ix29978 (.Y (nx29977), .A0 (label_6_output[9]), .A1 (
          booth_booth_integration_output_5_9), .B0 (nx11986), .B1 (nx13287)) ;
    dffr labelsregfile_label6_loop1_9_fx_reg_q (.Q (label_6_output[9]), .QB (
         \$dummy [354]), .D (nx21213), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_9 (.Q (label_6_input_9), .D (nx12000), .CLK (nx34523
          )) ;
    dffr reg_label_6_input_state_machine_9 (.Q (label_6_input_state_machine_9), 
         .QB (\$dummy [355]), .D (nx21203), .CLK (clk), .R (rst)) ;
    xnor2 ix11997 (.Y (nx11996), .A0 (nx11986), .A1 (nx30093)) ;
    oai22 ix11987 (.Y (nx11986), .A0 (nx29988), .A1 (nx30082), .B0 (nx30092), .B1 (
          nx29929)) ;
    aoi22 ix29989 (.Y (nx29988), .A0 (label_6_output[7]), .A1 (
          booth_booth_integration_output_5_7), .B0 (nx11922), .B1 (nx13285)) ;
    dffr labelsregfile_label6_loop1_7_fx_reg_q (.Q (label_6_output[7]), .QB (
         \$dummy [356]), .D (nx21173), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_7 (.Q (label_6_input_7), .D (nx11936), .CLK (nx34523
          )) ;
    dffr reg_label_6_input_state_machine_7 (.Q (label_6_input_state_machine_7), 
         .QB (\$dummy [357]), .D (nx21163), .CLK (clk), .R (rst)) ;
    xnor2 ix11933 (.Y (nx11932), .A0 (nx11922), .A1 (nx30078)) ;
    oai22 ix11923 (.Y (nx11922), .A0 (nx29999), .A1 (nx30067), .B0 (nx30077), .B1 (
          nx29931)) ;
    aoi22 ix30000 (.Y (nx29999), .A0 (label_6_output[5]), .A1 (
          booth_booth_integration_output_5_5), .B0 (nx11858), .B1 (nx13283)) ;
    dffr labelsregfile_label6_loop1_5_fx_reg_q (.Q (label_6_output[5]), .QB (
         \$dummy [358]), .D (nx21133), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_5 (.Q (label_6_input_5), .D (nx11872), .CLK (nx34521
          )) ;
    dffr reg_label_6_input_state_machine_5 (.Q (label_6_input_state_machine_5), 
         .QB (\$dummy [359]), .D (nx21123), .CLK (clk), .R (rst)) ;
    xnor2 ix11869 (.Y (nx11868), .A0 (nx11858), .A1 (nx30063)) ;
    oai22 ix11859 (.Y (nx11858), .A0 (nx30010), .A1 (nx30052), .B0 (nx30062), .B1 (
          nx29933)) ;
    aoi22 ix30011 (.Y (nx30010), .A0 (label_6_output[3]), .A1 (
          booth_booth_integration_output_5_3), .B0 (nx11794), .B1 (nx13279)) ;
    dffr labelsregfile_label6_loop1_3_fx_reg_q (.Q (label_6_output[3]), .QB (
         \$dummy [360]), .D (nx21093), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_3 (.Q (label_6_input_3), .D (nx11808), .CLK (nx34521
          )) ;
    dffr reg_label_6_input_state_machine_3 (.Q (label_6_input_state_machine_3), 
         .QB (\$dummy [361]), .D (nx21083), .CLK (clk), .R (rst)) ;
    xnor2 ix11805 (.Y (nx11804), .A0 (nx11794), .A1 (nx30048)) ;
    oai22 ix11795 (.Y (nx11794), .A0 (nx30021), .A1 (nx30037), .B0 (nx30047), .B1 (
          nx29935)) ;
    aoi32 ix30022 (.Y (nx30021), .A0 (label_6_output[0]), .A1 (nx35767), .A2 (
          nx13276), .B0 (label_6_output[1]), .B1 (
          booth_booth_integration_output_5_1)) ;
    dffr labelsregfile_label6_loop1_1_fx_reg_q (.Q (label_6_output[1]), .QB (
         \$dummy [362]), .D (nx21053), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_1 (.Q (label_6_input_1), .D (nx11744), .CLK (nx34521
          )) ;
    dffr reg_label_6_input_state_machine_1 (.Q (label_6_input_state_machine_1), 
         .QB (\$dummy [363]), .D (nx21043), .CLK (clk), .R (rst)) ;
    xor2 ix11741 (.Y (nx11740), .A0 (nx30032), .A1 (nx30034)) ;
    nand02 ix30033 (.Y (nx30032), .A0 (label_6_output[0]), .A1 (nx35767)) ;
    xnor2 ix30035 (.Y (nx30034), .A0 (booth_booth_integration_output_5_1), .A1 (
          label_6_output[1])) ;
    dffr labelsregfile_label6_loop1_2_fx_reg_q (.Q (label_6_output[2]), .QB (
         nx30047), .D (nx21073), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_2 (.Q (label_6_input_2), .D (nx11776), .CLK (nx34521
          )) ;
    dffr reg_label_6_input_state_machine_2 (.Q (label_6_input_state_machine_2), 
         .QB (\$dummy [364]), .D (nx21063), .CLK (clk), .R (rst)) ;
    xor2 ix11773 (.Y (nx11772), .A0 (nx30021), .A1 (nx30037)) ;
    xnor2 ix30049 (.Y (nx30048), .A0 (booth_booth_integration_output_5_3), .A1 (
          label_6_output[3])) ;
    dffr labelsregfile_label6_loop1_4_fx_reg_q (.Q (label_6_output[4]), .QB (
         nx30062), .D (nx21113), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_4 (.Q (label_6_input_4), .D (nx11840), .CLK (nx34521
          )) ;
    dffr reg_label_6_input_state_machine_4 (.Q (label_6_input_state_machine_4), 
         .QB (\$dummy [365]), .D (nx21103), .CLK (clk), .R (rst)) ;
    xor2 ix11837 (.Y (nx11836), .A0 (nx30010), .A1 (nx30052)) ;
    xnor2 ix30064 (.Y (nx30063), .A0 (booth_booth_integration_output_5_5), .A1 (
          label_6_output[5])) ;
    dffr labelsregfile_label6_loop1_6_fx_reg_q (.Q (label_6_output[6]), .QB (
         nx30077), .D (nx21153), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_6 (.Q (label_6_input_6), .D (nx11904), .CLK (nx34523
          )) ;
    dffr reg_label_6_input_state_machine_6 (.Q (label_6_input_state_machine_6), 
         .QB (\$dummy [366]), .D (nx21143), .CLK (clk), .R (rst)) ;
    xor2 ix11901 (.Y (nx11900), .A0 (nx29999), .A1 (nx30067)) ;
    xnor2 ix30079 (.Y (nx30078), .A0 (booth_booth_integration_output_5_7), .A1 (
          label_6_output[7])) ;
    dffr labelsregfile_label6_loop1_8_fx_reg_q (.Q (label_6_output[8]), .QB (
         nx30092), .D (nx21193), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_8 (.Q (label_6_input_8), .D (nx11968), .CLK (nx34523
          )) ;
    dffr reg_label_6_input_state_machine_8 (.Q (label_6_input_state_machine_8), 
         .QB (\$dummy [367]), .D (nx21183), .CLK (clk), .R (rst)) ;
    xor2 ix11965 (.Y (nx11964), .A0 (nx29988), .A1 (nx30082)) ;
    xnor2 ix30094 (.Y (nx30093), .A0 (booth_booth_integration_output_5_9), .A1 (
          label_6_output[9])) ;
    dffr labelsregfile_label6_loop1_10_fx_reg_q (.Q (label_6_output[10]), .QB (
         nx30107), .D (nx21233), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_10 (.Q (label_6_input_10), .D (nx12032), .CLK (
          nx34523)) ;
    dffr reg_label_6_input_state_machine_10 (.Q (label_6_input_state_machine_10)
         , .QB (\$dummy [368]), .D (nx21223), .CLK (clk), .R (rst)) ;
    xor2 ix12029 (.Y (nx12028), .A0 (nx29977), .A1 (nx30097)) ;
    xnor2 ix30109 (.Y (nx30108), .A0 (booth_booth_integration_output_5_11), .A1 (
          label_6_output[11])) ;
    dffr labelsregfile_label6_loop1_12_fx_reg_q (.Q (label_6_output[12]), .QB (
         nx30122), .D (nx21273), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_12 (.Q (label_6_input_12), .D (nx12096), .CLK (
          nx34523)) ;
    dffr reg_label_6_input_state_machine_12 (.Q (label_6_input_state_machine_12)
         , .QB (\$dummy [369]), .D (nx21263), .CLK (clk), .R (rst)) ;
    xor2 ix12093 (.Y (nx12092), .A0 (nx29966), .A1 (nx30112)) ;
    xnor2 ix30124 (.Y (nx30123), .A0 (booth_booth_integration_output_5_13), .A1 (
          label_6_output[13])) ;
    oai21 ix20474 (.Y (nx20473), .A0 (nx30132), .A1 (nx34767), .B0 (nx30134)) ;
    dff max_calc_reg_comparator_third_inp1_14 (.Q (
        max_calc_comparator_third_inp1_14), .QB (nx30132), .D (nx20473), .CLK (
        clk)) ;
    dffr labelsregfile_label5_loop1_14_fx_reg_q (.Q (label_5_output[14]), .QB (
         nx30318), .D (nx20463), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_14 (.Q (label_5_input_14), .D (nx10832), .CLK (
          nx34529)) ;
    dffr reg_label_5_input_state_machine_14 (.Q (label_5_input_state_machine_14)
         , .QB (\$dummy [370]), .D (nx19643), .CLK (clk), .R (rst)) ;
    xor2 ix10829 (.Y (nx10828), .A0 (nx30144), .A1 (nx30316)) ;
    aoi22 ix30145 (.Y (nx30144), .A0 (label_5_output[13]), .A1 (
          booth_booth_integration_output_4_13), .B0 (nx10792), .B1 (nx13253)) ;
    dffr labelsregfile_label5_loop1_13_fx_reg_q (.Q (label_5_output[13]), .QB (
         \$dummy [371]), .D (nx20453), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_13 (.Q (label_5_input_13), .D (nx10806), .CLK (
          nx34529)) ;
    dffr reg_label_5_input_state_machine_13 (.Q (label_5_input_state_machine_13)
         , .QB (\$dummy [372]), .D (nx20443), .CLK (clk), .R (rst)) ;
    xnor2 ix10803 (.Y (nx10802), .A0 (nx10792), .A1 (nx30312)) ;
    oai22 ix10793 (.Y (nx10792), .A0 (nx30155), .A1 (nx30301), .B0 (nx30311), .B1 (
          nx29484)) ;
    aoi22 ix30156 (.Y (nx30155), .A0 (label_5_output[11]), .A1 (
          booth_booth_integration_output_4_11), .B0 (nx10728), .B1 (nx13251)) ;
    dffr labelsregfile_label5_loop1_11_fx_reg_q (.Q (label_5_output[11]), .QB (
         \$dummy [373]), .D (nx20413), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_11 (.Q (label_5_input_11), .D (nx10742), .CLK (
          nx34527)) ;
    dffr reg_label_5_input_state_machine_11 (.Q (label_5_input_state_machine_11)
         , .QB (\$dummy [374]), .D (nx20403), .CLK (clk), .R (rst)) ;
    xnor2 ix10739 (.Y (nx10738), .A0 (nx10728), .A1 (nx30297)) ;
    oai22 ix10729 (.Y (nx10728), .A0 (nx30166), .A1 (nx30286), .B0 (nx30296), .B1 (
          nx29486)) ;
    aoi22 ix30167 (.Y (nx30166), .A0 (label_5_output[9]), .A1 (
          booth_booth_integration_output_4_9), .B0 (nx10664), .B1 (nx13249)) ;
    dffr labelsregfile_label5_loop1_9_fx_reg_q (.Q (label_5_output[9]), .QB (
         \$dummy [375]), .D (nx20373), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_9 (.Q (label_5_input_9), .D (nx10678), .CLK (nx34527
          )) ;
    dffr reg_label_5_input_state_machine_9 (.Q (label_5_input_state_machine_9), 
         .QB (\$dummy [376]), .D (nx20363), .CLK (clk), .R (rst)) ;
    xnor2 ix10675 (.Y (nx10674), .A0 (nx10664), .A1 (nx30282)) ;
    oai22 ix10665 (.Y (nx10664), .A0 (nx30177), .A1 (nx30271), .B0 (nx30281), .B1 (
          nx29488)) ;
    aoi22 ix30178 (.Y (nx30177), .A0 (label_5_output[7]), .A1 (
          booth_booth_integration_output_4_7), .B0 (nx10600), .B1 (nx13247)) ;
    dffr labelsregfile_label5_loop1_7_fx_reg_q (.Q (label_5_output[7]), .QB (
         \$dummy [377]), .D (nx20333), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_7 (.Q (label_5_input_7), .D (nx10614), .CLK (nx34527
          )) ;
    dffr reg_label_5_input_state_machine_7 (.Q (label_5_input_state_machine_7), 
         .QB (\$dummy [378]), .D (nx20323), .CLK (clk), .R (rst)) ;
    xnor2 ix10611 (.Y (nx10610), .A0 (nx10600), .A1 (nx30267)) ;
    oai22 ix10601 (.Y (nx10600), .A0 (nx30188), .A1 (nx30256), .B0 (nx30266), .B1 (
          nx29490)) ;
    aoi22 ix30189 (.Y (nx30188), .A0 (label_5_output[5]), .A1 (
          booth_booth_integration_output_4_5), .B0 (nx10536), .B1 (nx13243)) ;
    dffr labelsregfile_label5_loop1_5_fx_reg_q (.Q (label_5_output[5]), .QB (
         \$dummy [379]), .D (nx20293), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_5 (.Q (label_5_input_5), .D (nx10550), .CLK (nx34525
          )) ;
    dffr reg_label_5_input_state_machine_5 (.Q (label_5_input_state_machine_5), 
         .QB (\$dummy [380]), .D (nx20283), .CLK (clk), .R (rst)) ;
    xnor2 ix10547 (.Y (nx10546), .A0 (nx10536), .A1 (nx30252)) ;
    oai22 ix10537 (.Y (nx10536), .A0 (nx30199), .A1 (nx30241), .B0 (nx30251), .B1 (
          nx29492)) ;
    aoi22 ix30200 (.Y (nx30199), .A0 (label_5_output[3]), .A1 (
          booth_booth_integration_output_4_3), .B0 (nx10472), .B1 (nx13240)) ;
    dffr labelsregfile_label5_loop1_3_fx_reg_q (.Q (label_5_output[3]), .QB (
         \$dummy [381]), .D (nx20253), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_3 (.Q (label_5_input_3), .D (nx10486), .CLK (nx34525
          )) ;
    dffr reg_label_5_input_state_machine_3 (.Q (label_5_input_state_machine_3), 
         .QB (\$dummy [382]), .D (nx20243), .CLK (clk), .R (rst)) ;
    xnor2 ix10483 (.Y (nx10482), .A0 (nx10472), .A1 (nx30237)) ;
    oai22 ix10473 (.Y (nx10472), .A0 (nx30210), .A1 (nx30226), .B0 (nx30236), .B1 (
          nx29494)) ;
    aoi32 ix30211 (.Y (nx30210), .A0 (label_5_output[0]), .A1 (nx35763), .A2 (
          nx13238), .B0 (label_5_output[1]), .B1 (
          booth_booth_integration_output_4_1)) ;
    dffr labelsregfile_label5_loop1_1_fx_reg_q (.Q (label_5_output[1]), .QB (
         \$dummy [383]), .D (nx20213), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_1 (.Q (label_5_input_1), .D (nx10422), .CLK (nx34525
          )) ;
    dffr reg_label_5_input_state_machine_1 (.Q (label_5_input_state_machine_1), 
         .QB (\$dummy [384]), .D (nx20203), .CLK (clk), .R (rst)) ;
    xor2 ix10419 (.Y (nx10418), .A0 (nx30221), .A1 (nx30223)) ;
    nand02 ix30222 (.Y (nx30221), .A0 (label_5_output[0]), .A1 (nx35763)) ;
    xnor2 ix30224 (.Y (nx30223), .A0 (booth_booth_integration_output_4_1), .A1 (
          label_5_output[1])) ;
    dffr labelsregfile_label5_loop1_2_fx_reg_q (.Q (label_5_output[2]), .QB (
         nx30236), .D (nx20233), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_2 (.Q (label_5_input_2), .D (nx10454), .CLK (nx34525
          )) ;
    dffr reg_label_5_input_state_machine_2 (.Q (label_5_input_state_machine_2), 
         .QB (\$dummy [385]), .D (nx20223), .CLK (clk), .R (rst)) ;
    xor2 ix10451 (.Y (nx10450), .A0 (nx30210), .A1 (nx30226)) ;
    xnor2 ix30238 (.Y (nx30237), .A0 (booth_booth_integration_output_4_3), .A1 (
          label_5_output[3])) ;
    dffr labelsregfile_label5_loop1_4_fx_reg_q (.Q (label_5_output[4]), .QB (
         nx30251), .D (nx20273), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_4 (.Q (label_5_input_4), .D (nx10518), .CLK (nx34525
          )) ;
    dffr reg_label_5_input_state_machine_4 (.Q (label_5_input_state_machine_4), 
         .QB (\$dummy [386]), .D (nx20263), .CLK (clk), .R (rst)) ;
    xor2 ix10515 (.Y (nx10514), .A0 (nx30199), .A1 (nx30241)) ;
    xnor2 ix30253 (.Y (nx30252), .A0 (booth_booth_integration_output_4_5), .A1 (
          label_5_output[5])) ;
    dffr labelsregfile_label5_loop1_6_fx_reg_q (.Q (label_5_output[6]), .QB (
         nx30266), .D (nx20313), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_6 (.Q (label_5_input_6), .D (nx10582), .CLK (nx34527
          )) ;
    dffr reg_label_5_input_state_machine_6 (.Q (label_5_input_state_machine_6), 
         .QB (\$dummy [387]), .D (nx20303), .CLK (clk), .R (rst)) ;
    xor2 ix10579 (.Y (nx10578), .A0 (nx30188), .A1 (nx30256)) ;
    xnor2 ix30268 (.Y (nx30267), .A0 (booth_booth_integration_output_4_7), .A1 (
          label_5_output[7])) ;
    dffr labelsregfile_label5_loop1_8_fx_reg_q (.Q (label_5_output[8]), .QB (
         nx30281), .D (nx20353), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_8 (.Q (label_5_input_8), .D (nx10646), .CLK (nx34527
          )) ;
    dffr reg_label_5_input_state_machine_8 (.Q (label_5_input_state_machine_8), 
         .QB (\$dummy [388]), .D (nx20343), .CLK (clk), .R (rst)) ;
    xor2 ix10643 (.Y (nx10642), .A0 (nx30177), .A1 (nx30271)) ;
    xnor2 ix30283 (.Y (nx30282), .A0 (booth_booth_integration_output_4_9), .A1 (
          label_5_output[9])) ;
    dffr labelsregfile_label5_loop1_10_fx_reg_q (.Q (label_5_output[10]), .QB (
         nx30296), .D (nx20393), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_10 (.Q (label_5_input_10), .D (nx10710), .CLK (
          nx34527)) ;
    dffr reg_label_5_input_state_machine_10 (.Q (label_5_input_state_machine_10)
         , .QB (\$dummy [389]), .D (nx20383), .CLK (clk), .R (rst)) ;
    xor2 ix10707 (.Y (nx10706), .A0 (nx30166), .A1 (nx30286)) ;
    xnor2 ix30298 (.Y (nx30297), .A0 (booth_booth_integration_output_4_11), .A1 (
          label_5_output[11])) ;
    dffr labelsregfile_label5_loop1_12_fx_reg_q (.Q (label_5_output[12]), .QB (
         nx30311), .D (nx20433), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_12 (.Q (label_5_input_12), .D (nx10774), .CLK (
          nx34527)) ;
    dffr reg_label_5_input_state_machine_12 (.Q (label_5_input_state_machine_12)
         , .QB (\$dummy [390]), .D (nx20423), .CLK (clk), .R (rst)) ;
    xor2 ix10771 (.Y (nx10770), .A0 (nx30155), .A1 (nx30301)) ;
    xnor2 ix30313 (.Y (nx30312), .A0 (booth_booth_integration_output_4_13), .A1 (
          label_5_output[13])) ;
    oai22 ix12595 (.Y (nx12594), .A0 (nx30321), .A1 (nx30334), .B0 (
          max_calc_comparator_third_inp2_13), .B1 (nx30329)) ;
    oai21 ix21324 (.Y (nx21323), .A0 (nx30325), .A1 (nx34767), .B0 (nx30327)) ;
    dff max_calc_reg_comparator_third_inp2_13 (.Q (
        max_calc_comparator_third_inp2_13), .QB (nx30325), .D (nx21323), .CLK (
        clk)) ;
    nand03 ix30328 (.Y (nx30327), .A0 (label_6_output[13]), .A1 (nx35453), .A2 (
           nx34767)) ;
    dff max_calc_reg_comparator_third_inp1_13 (.Q (
        max_calc_comparator_third_inp1_13), .QB (nx30329), .D (nx21333), .CLK (
        clk)) ;
    oai21 ix21334 (.Y (nx21333), .A0 (nx30329), .A1 (nx34767), .B0 (nx30332)) ;
    nand03 ix30333 (.Y (nx30332), .A0 (label_5_output[13]), .A1 (nx35453), .A2 (
           nx34767)) ;
    aoi22 ix30335 (.Y (nx30334), .A0 (nx30336), .A1 (
          max_calc_comparator_third_inp1_12), .B0 (nx12220), .B1 (nx12578)) ;
    dff max_calc_reg_comparator_third_inp2_12 (.Q (\$dummy [391]), .QB (nx30336)
        , .D (nx21343), .CLK (clk)) ;
    oai21 ix21344 (.Y (nx21343), .A0 (nx30336), .A1 (nx34769), .B0 (nx30339)) ;
    oai21 ix21354 (.Y (nx21353), .A0 (nx30343), .A1 (nx34769), .B0 (nx30345)) ;
    dff max_calc_reg_comparator_third_inp1_12 (.Q (
        max_calc_comparator_third_inp1_12), .QB (nx30343), .D (nx21353), .CLK (
        clk)) ;
    oai22 ix12579 (.Y (nx12578), .A0 (nx30349), .A1 (nx30362), .B0 (
          max_calc_comparator_third_inp2_11), .B1 (nx30357)) ;
    oai21 ix21364 (.Y (nx21363), .A0 (nx30353), .A1 (nx34769), .B0 (nx30355)) ;
    dff max_calc_reg_comparator_third_inp2_11 (.Q (
        max_calc_comparator_third_inp2_11), .QB (nx30353), .D (nx21363), .CLK (
        clk)) ;
    nand03 ix30356 (.Y (nx30355), .A0 (label_6_output[11]), .A1 (nx35455), .A2 (
           nx34769)) ;
    dff max_calc_reg_comparator_third_inp1_11 (.Q (
        max_calc_comparator_third_inp1_11), .QB (nx30357), .D (nx21373), .CLK (
        clk)) ;
    oai21 ix21374 (.Y (nx21373), .A0 (nx30357), .A1 (nx34769), .B0 (nx30360)) ;
    nand03 ix30361 (.Y (nx30360), .A0 (label_5_output[11]), .A1 (nx35455), .A2 (
           nx34771)) ;
    aoi22 ix30363 (.Y (nx30362), .A0 (nx30364), .A1 (
          max_calc_comparator_third_inp1_10), .B0 (nx12264), .B1 (nx12562)) ;
    dff max_calc_reg_comparator_third_inp2_10 (.Q (\$dummy [392]), .QB (nx30364)
        , .D (nx21383), .CLK (clk)) ;
    oai21 ix21384 (.Y (nx21383), .A0 (nx30364), .A1 (nx34771), .B0 (nx30367)) ;
    oai21 ix21394 (.Y (nx21393), .A0 (nx30371), .A1 (nx34771), .B0 (nx30373)) ;
    dff max_calc_reg_comparator_third_inp1_10 (.Q (
        max_calc_comparator_third_inp1_10), .QB (nx30371), .D (nx21393), .CLK (
        clk)) ;
    oai22 ix12563 (.Y (nx12562), .A0 (nx30377), .A1 (nx30390), .B0 (
          max_calc_comparator_third_inp2_9), .B1 (nx30385)) ;
    oai21 ix21404 (.Y (nx21403), .A0 (nx30381), .A1 (nx34771), .B0 (nx30383)) ;
    dff max_calc_reg_comparator_third_inp2_9 (.Q (
        max_calc_comparator_third_inp2_9), .QB (nx30381), .D (nx21403), .CLK (
        clk)) ;
    nand03 ix30384 (.Y (nx30383), .A0 (label_6_output[9]), .A1 (nx35455), .A2 (
           nx34771)) ;
    dff max_calc_reg_comparator_third_inp1_9 (.Q (
        max_calc_comparator_third_inp1_9), .QB (nx30385), .D (nx21413), .CLK (
        clk)) ;
    oai21 ix21414 (.Y (nx21413), .A0 (nx30385), .A1 (nx34773), .B0 (nx30388)) ;
    nand03 ix30389 (.Y (nx30388), .A0 (label_5_output[9]), .A1 (nx35455), .A2 (
           nx34773)) ;
    aoi22 ix30391 (.Y (nx30390), .A0 (nx30392), .A1 (
          max_calc_comparator_third_inp1_8), .B0 (nx12308), .B1 (nx12546)) ;
    dff max_calc_reg_comparator_third_inp2_8 (.Q (\$dummy [393]), .QB (nx30392)
        , .D (nx21423), .CLK (clk)) ;
    oai21 ix21424 (.Y (nx21423), .A0 (nx30392), .A1 (nx34773), .B0 (nx30395)) ;
    oai21 ix21434 (.Y (nx21433), .A0 (nx30399), .A1 (nx34773), .B0 (nx30401)) ;
    dff max_calc_reg_comparator_third_inp1_8 (.Q (
        max_calc_comparator_third_inp1_8), .QB (nx30399), .D (nx21433), .CLK (
        clk)) ;
    oai22 ix12547 (.Y (nx12546), .A0 (nx30405), .A1 (nx30418), .B0 (
          max_calc_comparator_third_inp2_7), .B1 (nx30413)) ;
    oai21 ix21444 (.Y (nx21443), .A0 (nx30409), .A1 (nx34773), .B0 (nx30411)) ;
    dff max_calc_reg_comparator_third_inp2_7 (.Q (
        max_calc_comparator_third_inp2_7), .QB (nx30409), .D (nx21443), .CLK (
        clk)) ;
    nand03 ix30412 (.Y (nx30411), .A0 (label_6_output[7]), .A1 (nx35457), .A2 (
           nx34775)) ;
    dff max_calc_reg_comparator_third_inp1_7 (.Q (
        max_calc_comparator_third_inp1_7), .QB (nx30413), .D (nx21453), .CLK (
        clk)) ;
    oai21 ix21454 (.Y (nx21453), .A0 (nx30413), .A1 (nx34775), .B0 (nx30416)) ;
    nand03 ix30417 (.Y (nx30416), .A0 (label_5_output[7]), .A1 (nx35457), .A2 (
           nx34775)) ;
    aoi22 ix30419 (.Y (nx30418), .A0 (nx30420), .A1 (
          max_calc_comparator_third_inp1_6), .B0 (nx12352), .B1 (nx12530)) ;
    dff max_calc_reg_comparator_third_inp2_6 (.Q (\$dummy [394]), .QB (nx30420)
        , .D (nx21463), .CLK (clk)) ;
    oai21 ix21464 (.Y (nx21463), .A0 (nx30420), .A1 (nx34775), .B0 (nx30423)) ;
    oai21 ix21474 (.Y (nx21473), .A0 (nx30427), .A1 (nx34775), .B0 (nx30429)) ;
    dff max_calc_reg_comparator_third_inp1_6 (.Q (
        max_calc_comparator_third_inp1_6), .QB (nx30427), .D (nx21473), .CLK (
        clk)) ;
    oai22 ix12531 (.Y (nx12530), .A0 (nx30433), .A1 (nx30446), .B0 (
          max_calc_comparator_third_inp2_5), .B1 (nx30441)) ;
    oai21 ix21484 (.Y (nx21483), .A0 (nx30437), .A1 (nx34777), .B0 (nx30439)) ;
    dff max_calc_reg_comparator_third_inp2_5 (.Q (
        max_calc_comparator_third_inp2_5), .QB (nx30437), .D (nx21483), .CLK (
        clk)) ;
    nand03 ix30440 (.Y (nx30439), .A0 (label_6_output[5]), .A1 (nx35457), .A2 (
           nx34777)) ;
    dff max_calc_reg_comparator_third_inp1_5 (.Q (
        max_calc_comparator_third_inp1_5), .QB (nx30441), .D (nx21493), .CLK (
        clk)) ;
    oai21 ix21494 (.Y (nx21493), .A0 (nx30441), .A1 (nx34777), .B0 (nx30444)) ;
    nand03 ix30445 (.Y (nx30444), .A0 (label_5_output[5]), .A1 (nx35459), .A2 (
           nx34777)) ;
    aoi22 ix30447 (.Y (nx30446), .A0 (nx30448), .A1 (
          max_calc_comparator_third_inp1_4), .B0 (nx12396), .B1 (nx12514)) ;
    dff max_calc_reg_comparator_third_inp2_4 (.Q (\$dummy [395]), .QB (nx30448)
        , .D (nx21503), .CLK (clk)) ;
    oai21 ix21504 (.Y (nx21503), .A0 (nx30448), .A1 (nx34777), .B0 (nx30451)) ;
    oai21 ix21514 (.Y (nx21513), .A0 (nx30455), .A1 (nx34777), .B0 (nx30457)) ;
    dff max_calc_reg_comparator_third_inp1_4 (.Q (
        max_calc_comparator_third_inp1_4), .QB (nx30455), .D (nx21513), .CLK (
        clk)) ;
    oai22 ix12515 (.Y (nx12514), .A0 (nx30461), .A1 (nx30474), .B0 (
          max_calc_comparator_third_inp2_3), .B1 (nx30469)) ;
    oai21 ix21524 (.Y (nx21523), .A0 (nx30465), .A1 (nx34779), .B0 (nx30467)) ;
    dff max_calc_reg_comparator_third_inp2_3 (.Q (
        max_calc_comparator_third_inp2_3), .QB (nx30465), .D (nx21523), .CLK (
        clk)) ;
    nand03 ix30468 (.Y (nx30467), .A0 (label_6_output[3]), .A1 (nx35459), .A2 (
           nx34779)) ;
    dff max_calc_reg_comparator_third_inp1_3 (.Q (
        max_calc_comparator_third_inp1_3), .QB (nx30469), .D (nx21533), .CLK (
        clk)) ;
    oai21 ix21534 (.Y (nx21533), .A0 (nx30469), .A1 (nx34779), .B0 (nx30472)) ;
    nand03 ix30473 (.Y (nx30472), .A0 (label_5_output[3]), .A1 (nx35459), .A2 (
           nx34779)) ;
    aoi22 ix30475 (.Y (nx30474), .A0 (nx30476), .A1 (
          max_calc_comparator_third_inp1_2), .B0 (nx12440), .B1 (nx12498)) ;
    dff max_calc_reg_comparator_third_inp2_2 (.Q (\$dummy [396]), .QB (nx30476)
        , .D (nx21543), .CLK (clk)) ;
    oai21 ix21544 (.Y (nx21543), .A0 (nx30476), .A1 (nx34779), .B0 (nx30479)) ;
    oai21 ix21554 (.Y (nx21553), .A0 (nx30483), .A1 (nx34781), .B0 (nx30485)) ;
    dff max_calc_reg_comparator_third_inp1_2 (.Q (
        max_calc_comparator_third_inp1_2), .QB (nx30483), .D (nx21553), .CLK (
        clk)) ;
    oai21 ix12499 (.Y (nx12498), .A0 (max_calc_comparator_third_inp2_1), .A1 (
          nx30495), .B0 (nx30500)) ;
    oai21 ix21564 (.Y (nx21563), .A0 (nx30491), .A1 (nx34781), .B0 (nx30493)) ;
    dff max_calc_reg_comparator_third_inp2_1 (.Q (
        max_calc_comparator_third_inp2_1), .QB (nx30491), .D (nx21563), .CLK (
        clk)) ;
    nand03 ix30494 (.Y (nx30493), .A0 (label_6_output[1]), .A1 (nx35461), .A2 (
           nx34781)) ;
    dff max_calc_reg_comparator_third_inp1_1 (.Q (\$dummy [397]), .QB (nx30495)
        , .D (nx21573), .CLK (clk)) ;
    oai21 ix21574 (.Y (nx21573), .A0 (nx30495), .A1 (nx34781), .B0 (nx30498)) ;
    nand03 ix30499 (.Y (nx30498), .A0 (label_5_output[1]), .A1 (nx35461), .A2 (
           nx34781)) ;
    oai21 ix30501 (.Y (nx30500), .A0 (nx29502), .A1 (
          max_calc_comparator_third_inp1_0), .B0 (nx12462)) ;
    oai21 ix21624 (.Y (nx21623), .A0 (nx30506), .A1 (nx34781), .B0 (nx30508)) ;
    dff max_calc_reg_comparator_third_inp2_15 (.Q (\$dummy [398]), .QB (nx30506)
        , .D (nx21623), .CLK (clk)) ;
    nand03 ix30509 (.Y (nx30508), .A0 (label_6_output[15]), .A1 (nx35461), .A2 (
           nx34783)) ;
    dffr labelsregfile_label6_loop1_15_fx_reg_q (.Q (label_6_output[15]), .QB (
         \$dummy [399]), .D (nx21613), .CLK (clk), .R (rst)) ;
    latch lat_label_6_input_15 (.Q (label_6_input_15), .D (nx12624), .CLK (
          nx34529)) ;
    dffr reg_label_6_input_state_machine_15 (.Q (label_6_input_state_machine_15)
         , .QB (\$dummy [400]), .D (nx21603), .CLK (clk), .R (rst)) ;
    xnor2 ix12621 (.Y (nx12620), .A0 (nx12616), .A1 (nx30519)) ;
    oai22 ix12617 (.Y (nx12616), .A0 (nx29955), .A1 (nx30127), .B0 (nx30129), .B1 (
          nx29923)) ;
    oai21 ix21654 (.Y (nx21653), .A0 (nx30524), .A1 (nx34783), .B0 (nx30526)) ;
    dff max_calc_reg_comparator_third_inp1_15 (.Q (\$dummy [401]), .QB (nx30524)
        , .D (nx21653), .CLK (clk)) ;
    nand03 ix30527 (.Y (nx30526), .A0 (label_5_output[15]), .A1 (nx35461), .A2 (
           nx34783)) ;
    dffr labelsregfile_label5_loop1_15_fx_reg_q (.Q (label_5_output[15]), .QB (
         \$dummy [402]), .D (nx21643), .CLK (clk), .R (rst)) ;
    latch lat_label_5_input_15 (.Q (label_5_input_15), .D (nx12666), .CLK (
          nx34529)) ;
    dffr reg_label_5_input_state_machine_15 (.Q (label_5_input_state_machine_15)
         , .QB (\$dummy [403]), .D (nx21633), .CLK (clk), .R (rst)) ;
    xnor2 ix12663 (.Y (nx12662), .A0 (nx12658), .A1 (nx30537)) ;
    oai22 ix12659 (.Y (nx12658), .A0 (nx30144), .A1 (nx30316), .B0 (nx30318), .B1 (
          nx29482)) ;
    dff max_calc_reg_ans3_0 (.Q (max_calc_ans3_0), .QB (\$dummy [404]), .D (
        nx24263), .CLK (clk)) ;
    oai21 ix24254 (.Y (nx24253), .A0 (nx30546), .A1 (nx34783), .B0 (nx30548)) ;
    dff max_calc_reg_comparator_second_inp2_0 (.Q (\$dummy [405]), .QB (nx30546)
        , .D (nx24253), .CLK (clk)) ;
    nand03 ix30549 (.Y (nx30548), .A0 (nx35175), .A1 (nx16896), .A2 (nx34801)) ;
    dffr labelsregfile_label4_loop1_0_fx_reg_q (.Q (label_4_output[0]), .QB (
         \$dummy [406]), .D (nx14673), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_0 (.Q (label_4_input_0), .D (nx1744), .CLK (nx34529)
          ) ;
    oai21 ix1745 (.Y (nx1744), .A0 (nx30555), .A1 (nx34429), .B0 (nx30559)) ;
    dffr reg_label_4_input_state_machine_0 (.Q (label_4_input_state_machine_0), 
         .QB (nx30555), .D (nx14663), .CLK (clk), .R (rst)) ;
    oai21 ix30560 (.Y (nx30559), .A0 (nx35719), .A1 (label_4_output[0]), .B0 (
          nx1732)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_3_1), .QB (\$dummy [407]), .D (nx14643)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_3_2), .QB (nx30980), .D (nx14633), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_3_3), .QB (\$dummy [408]), .D (nx14623)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_3_4), .QB (nx30978), .D (nx14613), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_3_5), .QB (\$dummy [409]), .D (nx14603)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_3_6), .QB (nx30976), .D (nx14593), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_3_7), .QB (\$dummy [410]), .D (nx14583)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_3_8), .QB (nx30974), .D (nx14573), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_3_9), .QB (\$dummy [411]), .D (nx14563)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_3_10), .QB (nx30972), .D (nx14553), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_3_11), .QB (\$dummy [412]), .D (nx14543)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_3_12), .QB (nx30970), .D (nx14533), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_3_13), .QB (\$dummy [413]), .D (nx14523)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_3_14), .QB (nx30968), .D (nx14513), .CLK (
         clk), .R (rst)) ;
    aoi22 ix30609 (.Y (nx30608), .A0 (mdr_data_out[15]), .A1 (nx34571), .B0 (
          nx1530), .B1 (nx1536)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_reg_output_0), .QB (\$dummy [414]), .D (
         nx14153), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_3_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_3_shift_Reg_count_0), .QB (\$dummy [415]), .D (
            nx14139), .CLK (clk), .S (nx34487)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_reg_output_9), .QB (\$dummy [416]), .D (
         nx14333), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_9), .QB (\$dummy [417]), .D (
         nx14323), .CLK (clk), .R (nx34487)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_8), .QB (\$dummy [418]), .D (
         nx14313), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_8), .QB (\$dummy [419]), .D (
         nx14303), .CLK (clk), .R (nx34487)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_7), .QB (\$dummy [420]), .D (
         nx14293), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_7), .QB (\$dummy [421]), .D (
         nx14283), .CLK (clk), .R (nx34485)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_6), .QB (\$dummy [422]), .D (
         nx14273), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_6), .QB (\$dummy [423]), .D (
         nx14263), .CLK (clk), .R (nx34485)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_5), .QB (\$dummy [424]), .D (
         nx14253), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_5), .QB (\$dummy [425]), .D (
         nx14243), .CLK (clk), .R (nx34485)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_4), .QB (\$dummy [426]), .D (
         nx14233), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_4), .QB (\$dummy [427]), .D (
         nx14223), .CLK (clk), .R (nx34485)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_3), .QB (\$dummy [428]), .D (
         nx14213), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_3), .QB (\$dummy [429]), .D (
         nx14203), .CLK (clk), .R (nx34485)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_2), .QB (\$dummy [430]), .D (
         nx14193), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_2), .QB (\$dummy [431]), .D (
         nx14183), .CLK (clk), .R (nx34485)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_3_shift_Reg_output_1), .QB (\$dummy [432]), .D (
         nx14173), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_3_shift_Reg_count_1), .QB (\$dummy [433]), .D (
         nx14163), .CLK (clk), .R (nx34483)) ;
    nand02 ix14134 (.Y (nx14133), .A0 (nx35831), .A1 (nx34557)) ;
    dffs_ni booth_booth_integrtaion_3_shift_Reg_reg_en (.Q (\$dummy [434]), .QB (
            nx30655), .D (nx14133), .CLK (clk), .S (nx34485)) ;
    nand02 ix1531 (.Y (nx1530), .A0 (nx30676), .A1 (nx30688)) ;
    oai21 ix30677 (.Y (nx30676), .A0 (nx34585), .A1 (nx34579), .B0 (
          mdr_data_out[64])) ;
    oai21 ix14344 (.Y (nx14343), .A0 (nx30681), .A1 (nx35499), .B0 (nx30683)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [435]), .QB (
         nx30681), .D (nx14343), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [436]), .QB (
         nx30685), .D (nx14653), .CLK (clk), .R (rst)) ;
    xnor2 ix30693 (.Y (nx30692), .A0 (nx1000), .A1 (nx12913)) ;
    oai21 ix14484 (.Y (nx14483), .A0 (nx30698), .A1 (nx35499), .B0 (nx30700)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_17), .QB (nx30698), .D (nx14483)
         , .CLK (clk), .R (rst)) ;
    nand03 ix30701 (.Y (nx30700), .A0 (nx35507), .A1 (nx1508), .A2 (nx36147)) ;
    xnor2 ix1509 (.Y (nx1508), .A0 (nx30703), .A1 (nx12915)) ;
    aoi22 ix30704 (.Y (nx30703), .A0 (booth_booth_integrtaion_3_booth_output_17)
          , .A1 (nx1024), .B0 (nx1000), .B1 (nx12913)) ;
    nand02 ix1009 (.Y (nx1008), .A0 (mdr_data_out[65]), .A1 (mdr_data_out[64])
           ) ;
    or02 ix30708 (.Y (nx30707), .A0 (mdr_data_out[64]), .A1 (mdr_data_out[65])
         ) ;
    xnor2 ix30714 (.Y (nx30713), .A0 (nx1052), .A1 (nx12917)) ;
    oai22 ix1053 (.Y (nx1052), .A0 (nx30703), .A1 (nx30716), .B0 (nx30723), .B1 (
          nx35511)) ;
    aoi32 ix30719 (.Y (nx30718), .A0 (nx1034), .A1 (nx34585), .A2 (nx30721), .B0 (
          mdr_data_out[66]), .B1 (nx34579)) ;
    oai21 ix1035 (.Y (nx1034), .A0 (mdr_data_out[64]), .A1 (mdr_data_out[65]), .B0 (
          mdr_data_out[66])) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_18), .QB (nx30723), .D (nx14473)
         , .CLK (clk), .R (rst)) ;
    oai21 ix14464 (.Y (nx14463), .A0 (nx30728), .A1 (nx35499), .B0 (nx30730)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_19), .QB (nx30728), .D (nx14463)
         , .CLK (clk), .R (rst)) ;
    nand03 ix30731 (.Y (nx30730), .A0 (nx35507), .A1 (nx1484), .A2 (nx36147)) ;
    xnor2 ix1485 (.Y (nx1484), .A0 (nx30733), .A1 (nx12919)) ;
    aoi22 ix30734 (.Y (nx30733), .A0 (booth_booth_integrtaion_3_booth_output_19)
          , .A1 (nx1072), .B0 (nx1052), .B1 (nx12917)) ;
    nor02ii ix30737 (.Y (nx30736), .A0 (nx1038), .A1 (mdr_data_out[67])) ;
    nor03_2x ix1039 (.Y (nx1038), .A0 (mdr_data_out[66]), .A1 (mdr_data_out[64])
             , .A2 (mdr_data_out[65])) ;
    nor04 ix1063 (.Y (nx1062), .A0 (mdr_data_out[67]), .A1 (mdr_data_out[66]), .A2 (
          mdr_data_out[64]), .A3 (mdr_data_out[65])) ;
    xnor2 ix30751 (.Y (nx30750), .A0 (nx1100), .A1 (nx12921)) ;
    oai22 ix1101 (.Y (nx1100), .A0 (nx30733), .A1 (nx30753), .B0 (nx30762), .B1 (
          nx35513)) ;
    aoi32 ix30756 (.Y (nx30755), .A0 (nx1082), .A1 (nx34585), .A2 (nx30760), .B0 (
          mdr_data_out[68]), .B1 (nx34579)) ;
    nand02 ix1083 (.Y (nx1082), .A0 (nx30758), .A1 (mdr_data_out[68])) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_20), .QB (nx30762), .D (nx14453)
         , .CLK (clk), .R (rst)) ;
    oai21 ix14444 (.Y (nx14443), .A0 (nx30767), .A1 (nx35499), .B0 (nx30769)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_21), .QB (nx30767), .D (nx14443)
         , .CLK (clk), .R (rst)) ;
    nand03 ix30770 (.Y (nx30769), .A0 (nx35507), .A1 (nx1460), .A2 (nx36147)) ;
    xnor2 ix1461 (.Y (nx1460), .A0 (nx30772), .A1 (nx12922)) ;
    aoi22 ix30773 (.Y (nx30772), .A0 (booth_booth_integrtaion_3_booth_output_21)
          , .A1 (nx1120), .B0 (nx1100), .B1 (nx12921)) ;
    nor02ii ix30776 (.Y (nx30775), .A0 (nx1086), .A1 (mdr_data_out[69])) ;
    nor02ii ix1087 (.Y (nx1086), .A0 (mdr_data_out[68]), .A1 (nx1062)) ;
    nor02ii ix1111 (.Y (nx1110), .A0 (mdr_data_out[69]), .A1 (nx1086)) ;
    xnor2 ix30786 (.Y (nx30785), .A0 (nx1148), .A1 (nx12923)) ;
    oai22 ix1149 (.Y (nx1148), .A0 (nx30772), .A1 (nx30788), .B0 (nx30797), .B1 (
          nx35515)) ;
    aoi32 ix30791 (.Y (nx30790), .A0 (nx1130), .A1 (nx34585), .A2 (nx30795), .B0 (
          mdr_data_out[70]), .B1 (nx34579)) ;
    nand02 ix1131 (.Y (nx1130), .A0 (nx30793), .A1 (mdr_data_out[70])) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_22), .QB (nx30797), .D (nx14433)
         , .CLK (clk), .R (rst)) ;
    oai21 ix14424 (.Y (nx14423), .A0 (nx30802), .A1 (nx35499), .B0 (nx30804)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_23), .QB (nx30802), .D (nx14423)
         , .CLK (clk), .R (rst)) ;
    nand03 ix30805 (.Y (nx30804), .A0 (nx35507), .A1 (nx1436), .A2 (nx35501)) ;
    xnor2 ix1437 (.Y (nx1436), .A0 (nx30807), .A1 (nx12925)) ;
    aoi22 ix30808 (.Y (nx30807), .A0 (booth_booth_integrtaion_3_booth_output_23)
          , .A1 (nx1168), .B0 (nx1148), .B1 (nx12923)) ;
    nor02ii ix30811 (.Y (nx30810), .A0 (nx1134), .A1 (mdr_data_out[71])) ;
    nor02ii ix1135 (.Y (nx1134), .A0 (mdr_data_out[70]), .A1 (nx1110)) ;
    nor02ii ix1159 (.Y (nx1158), .A0 (mdr_data_out[71]), .A1 (nx1134)) ;
    xnor2 ix30821 (.Y (nx30820), .A0 (nx1196), .A1 (nx12927)) ;
    oai22 ix1197 (.Y (nx1196), .A0 (nx30807), .A1 (nx30823), .B0 (nx30832), .B1 (
          nx35517)) ;
    aoi32 ix30826 (.Y (nx30825), .A0 (nx1178), .A1 (nx34585), .A2 (nx30830), .B0 (
          mdr_data_out[72]), .B1 (nx34579)) ;
    nand02 ix1179 (.Y (nx1178), .A0 (nx30828), .A1 (mdr_data_out[72])) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_24), .QB (nx30832), .D (nx14413)
         , .CLK (clk), .R (rst)) ;
    oai21 ix14404 (.Y (nx14403), .A0 (nx30837), .A1 (nx35501), .B0 (nx30839)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_25), .QB (nx30837), .D (nx14403)
         , .CLK (clk), .R (rst)) ;
    nand03 ix30840 (.Y (nx30839), .A0 (nx35507), .A1 (nx1412), .A2 (nx35501)) ;
    xnor2 ix1413 (.Y (nx1412), .A0 (nx30842), .A1 (nx12929)) ;
    aoi22 ix30843 (.Y (nx30842), .A0 (booth_booth_integrtaion_3_booth_output_25)
          , .A1 (nx1216), .B0 (nx1196), .B1 (nx12927)) ;
    nor02ii ix30846 (.Y (nx30845), .A0 (nx1182), .A1 (mdr_data_out[73])) ;
    nor02ii ix1183 (.Y (nx1182), .A0 (mdr_data_out[72]), .A1 (nx1158)) ;
    nor02ii ix1207 (.Y (nx1206), .A0 (mdr_data_out[73]), .A1 (nx1182)) ;
    xnor2 ix30856 (.Y (nx30855), .A0 (nx1244), .A1 (nx12930)) ;
    oai22 ix1245 (.Y (nx1244), .A0 (nx30842), .A1 (nx30858), .B0 (nx30867), .B1 (
          nx35519)) ;
    aoi32 ix30861 (.Y (nx30860), .A0 (nx1226), .A1 (nx34585), .A2 (nx30865), .B0 (
          mdr_data_out[74]), .B1 (nx34579)) ;
    nand02 ix1227 (.Y (nx1226), .A0 (nx30863), .A1 (mdr_data_out[74])) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_26), .QB (nx30867), .D (nx14393)
         , .CLK (clk), .R (rst)) ;
    oai21 ix14384 (.Y (nx14383), .A0 (nx30872), .A1 (nx35501), .B0 (nx30874)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_27), .QB (nx30872), .D (nx14383)
         , .CLK (clk), .R (rst)) ;
    nand03 ix30875 (.Y (nx30874), .A0 (nx35507), .A1 (nx1388), .A2 (nx35501)) ;
    xnor2 ix1389 (.Y (nx1388), .A0 (nx30877), .A1 (nx12931)) ;
    aoi22 ix30878 (.Y (nx30877), .A0 (booth_booth_integrtaion_3_booth_output_27)
          , .A1 (nx1264), .B0 (nx1244), .B1 (nx12930)) ;
    nor02ii ix30881 (.Y (nx30880), .A0 (nx1230), .A1 (mdr_data_out[75])) ;
    nor02ii ix1231 (.Y (nx1230), .A0 (mdr_data_out[74]), .A1 (nx1206)) ;
    nor02ii ix1255 (.Y (nx1254), .A0 (mdr_data_out[75]), .A1 (nx1230)) ;
    xnor2 ix30891 (.Y (nx30890), .A0 (nx1292), .A1 (nx12933)) ;
    oai22 ix1293 (.Y (nx1292), .A0 (nx30877), .A1 (nx30893), .B0 (nx30902), .B1 (
          nx35521)) ;
    aoi32 ix30896 (.Y (nx30895), .A0 (nx1274), .A1 (nx34585), .A2 (nx30900), .B0 (
          mdr_data_out[76]), .B1 (nx34579)) ;
    nand02 ix1275 (.Y (nx1274), .A0 (nx30898), .A1 (mdr_data_out[76])) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_28), .QB (nx30902), .D (nx14373)
         , .CLK (clk), .R (rst)) ;
    oai21 ix14364 (.Y (nx14363), .A0 (nx30907), .A1 (nx35501), .B0 (nx30909)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_29), .QB (nx30907), .D (nx14363)
         , .CLK (clk), .R (rst)) ;
    nand03 ix30910 (.Y (nx30909), .A0 (nx36155), .A1 (nx1364), .A2 (nx35501)) ;
    xnor2 ix1365 (.Y (nx1364), .A0 (nx30912), .A1 (nx12935)) ;
    aoi22 ix30913 (.Y (nx30912), .A0 (booth_booth_integrtaion_3_booth_output_29)
          , .A1 (nx1312), .B0 (nx1292), .B1 (nx12933)) ;
    nor02ii ix30916 (.Y (nx30915), .A0 (nx1278), .A1 (mdr_data_out[77])) ;
    nor02ii ix1279 (.Y (nx1278), .A0 (mdr_data_out[76]), .A1 (nx1254)) ;
    nor02ii ix1303 (.Y (nx1302), .A0 (mdr_data_out[77]), .A1 (nx1278)) ;
    xnor2 ix30926 (.Y (nx30925), .A0 (nx1340), .A1 (nx1350)) ;
    oai22 ix1341 (.Y (nx1340), .A0 (nx30912), .A1 (nx30928), .B0 (nx30937), .B1 (
          nx35523)) ;
    aoi32 ix30931 (.Y (nx30930), .A0 (nx1322), .A1 (nx34587), .A2 (nx30935), .B0 (
          mdr_data_out[78]), .B1 (nx34581)) ;
    nand02 ix1323 (.Y (nx1322), .A0 (nx30933), .A1 (mdr_data_out[78])) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_31), .QB (nx30937), .D (nx14353)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix30941 (.Y (nx30940), .A0 (mdr_data_out[79]), .A1 (nx34581), .B0 (
          nx34587), .B1 (nx1342)) ;
    xnor2 ix1343 (.Y (nx1342), .A0 (mdr_data_out[79]), .A1 (nx1326)) ;
    nor02ii ix1327 (.Y (nx1326), .A0 (mdr_data_out[78]), .A1 (nx1302)) ;
    aoi32 ix30945 (.Y (nx30944), .A0 (nx1298), .A1 (nx34587), .A2 (nx30933), .B0 (
          mdr_data_out[77]), .B1 (nx34581)) ;
    aoi32 ix30948 (.Y (nx30947), .A0 (nx1250), .A1 (nx34587), .A2 (nx30898), .B0 (
          mdr_data_out[75]), .B1 (nx34581)) ;
    aoi32 ix30951 (.Y (nx30950), .A0 (nx1202), .A1 (nx34587), .A2 (nx30863), .B0 (
          mdr_data_out[73]), .B1 (nx34581)) ;
    aoi32 ix30954 (.Y (nx30953), .A0 (nx1154), .A1 (nx34587), .A2 (nx30828), .B0 (
          mdr_data_out[71]), .B1 (nx34581)) ;
    aoi32 ix30957 (.Y (nx30956), .A0 (nx1106), .A1 (nx34587), .A2 (nx30793), .B0 (
          mdr_data_out[69]), .B1 (nx34581)) ;
    aoi32 ix30960 (.Y (nx30959), .A0 (nx1058), .A1 (nx994), .A2 (nx30758), .B0 (
          mdr_data_out[67]), .B1 (nx34583)) ;
    aoi32 ix30963 (.Y (nx30962), .A0 (nx1008), .A1 (nx994), .A2 (nx30707), .B0 (
          mdr_data_out[65]), .B1 (nx34583)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_3_booth_output_16), .QB (nx30688), .D (nx14493)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_3_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_3_15), .QB (nx30966), .D (nx14503), .CLK (
         clk), .R (rst)) ;
    aoi21 ix1733 (.Y (nx1732), .A0 (label_4_output[0]), .A1 (nx35719), .B0 (
          nx35919)) ;
    oai21 ix23634 (.Y (nx23633), .A0 (nx30990), .A1 (nx34783), .B0 (nx30992)) ;
    dff max_calc_reg_comparator_fourth_inp1_0 (.Q (
        max_calc_comparator_fourth_inp1_0), .QB (nx30990), .D (nx23633), .CLK (
        clk)) ;
    nand03 ix30993 (.Y (nx30992), .A0 (label_7_output[0]), .A1 (nx35461), .A2 (
           nx34783)) ;
    dffr labelsregfile_label7_loop1_0_fx_reg_q (.Q (label_7_output[0]), .QB (
         \$dummy [437]), .D (nx22233), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_0 (.Q (label_7_input_0), .D (nx13586), .CLK (nx34529
          )) ;
    oai21 ix13587 (.Y (nx13586), .A0 (nx30998), .A1 (nx34429), .B0 (nx31002)) ;
    dffr reg_label_7_input_state_machine_0 (.Q (label_7_input_state_machine_0), 
         .QB (nx30998), .D (nx22223), .CLK (clk), .R (rst)) ;
    oai21 ix31003 (.Y (nx31002), .A0 (nx35771), .A1 (label_7_output[0]), .B0 (
          nx13574)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_6_1), .QB (\$dummy [438]), .D (nx22203)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_6_2), .QB (nx31423), .D (nx22193), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_6_3), .QB (\$dummy [439]), .D (nx22183)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_6_4), .QB (nx31421), .D (nx22173), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_6_5), .QB (\$dummy [440]), .D (nx22163)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_6_6), .QB (nx31419), .D (nx22153), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_6_7), .QB (\$dummy [441]), .D (nx22143)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_6_8), .QB (nx31417), .D (nx22133), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_6_9), .QB (\$dummy [442]), .D (nx22123)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_6_10), .QB (nx31415), .D (nx22113), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_6_11), .QB (\$dummy [443]), .D (nx22103)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_6_12), .QB (nx31413), .D (nx22093), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_6_13), .QB (\$dummy [444]), .D (nx22083)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_6_14), .QB (nx31411), .D (nx22073), .CLK (
         clk), .R (rst)) ;
    aoi22 ix31052 (.Y (nx31051), .A0 (mdr_data_out[15]), .A1 (nx35011), .B0 (
          nx13372), .B1 (nx13378)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_reg_output_0), .QB (\$dummy [445]), .D (
         nx21713), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_6_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_6_shift_Reg_count_0), .QB (\$dummy [446]), .D (
            nx21699), .CLK (clk), .S (nx34489)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_reg_output_9), .QB (\$dummy [447]), .D (
         nx21893), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_9), .QB (\$dummy [448]), .D (
         nx21883), .CLK (clk), .R (nx34489)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_8), .QB (\$dummy [449]), .D (
         nx21873), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_8), .QB (\$dummy [450]), .D (
         nx21863), .CLK (clk), .R (nx34489)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_7), .QB (\$dummy [451]), .D (
         nx21853), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_7), .QB (\$dummy [452]), .D (
         nx21843), .CLK (clk), .R (nx34489)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_6), .QB (\$dummy [453]), .D (
         nx21833), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_6), .QB (\$dummy [454]), .D (
         nx21823), .CLK (clk), .R (nx34489)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_5), .QB (\$dummy [455]), .D (
         nx21813), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_5), .QB (\$dummy [456]), .D (
         nx21803), .CLK (clk), .R (nx34489)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_4), .QB (\$dummy [457]), .D (
         nx21793), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_4), .QB (\$dummy [458]), .D (
         nx21783), .CLK (clk), .R (nx34489)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_3), .QB (\$dummy [459]), .D (
         nx21773), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_3), .QB (\$dummy [460]), .D (
         nx21763), .CLK (clk), .R (nx34487)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_2), .QB (\$dummy [461]), .D (
         nx21753), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_2), .QB (\$dummy [462]), .D (
         nx21743), .CLK (clk), .R (nx34487)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_6_shift_Reg_output_1), .QB (\$dummy [463]), .D (
         nx21733), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_6_shift_Reg_count_1), .QB (\$dummy [464]), .D (
         nx21723), .CLK (clk), .R (nx34487)) ;
    nand02 ix21694 (.Y (nx21693), .A0 (nx35835), .A1 (nx34997)) ;
    dffs_ni booth_booth_integrtaion_6_shift_Reg_reg_en (.Q (\$dummy [465]), .QB (
            nx31098), .D (nx21693), .CLK (clk), .S (nx34487)) ;
    nand02 ix13373 (.Y (nx13372), .A0 (nx31119), .A1 (nx31131)) ;
    oai21 ix31120 (.Y (nx31119), .A0 (nx35025), .A1 (nx35019), .B0 (
          mdr_data_out[112])) ;
    oai21 ix21904 (.Y (nx21903), .A0 (nx31124), .A1 (nx35525), .B0 (nx31126)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [466]), .QB (
         nx31124), .D (nx21903), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [467]), .QB (
         nx31128), .D (nx22213), .CLK (clk), .R (rst)) ;
    xnor2 ix31136 (.Y (nx31135), .A0 (nx12842), .A1 (nx13296)) ;
    oai21 ix22044 (.Y (nx22043), .A0 (nx31141), .A1 (nx35525), .B0 (nx31143)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_17), .QB (nx31141), .D (nx22043)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31144 (.Y (nx31143), .A0 (nx35533), .A1 (nx13350), .A2 (nx36163)) ;
    xnor2 ix13351 (.Y (nx13350), .A0 (nx31146), .A1 (nx13297)) ;
    aoi22 ix31147 (.Y (nx31146), .A0 (booth_booth_integrtaion_6_booth_output_17)
          , .A1 (nx12866), .B0 (nx12842), .B1 (nx13296)) ;
    nand02 ix12851 (.Y (nx12850), .A0 (mdr_data_out[113]), .A1 (
           mdr_data_out[112])) ;
    or02 ix31151 (.Y (nx31150), .A0 (mdr_data_out[112]), .A1 (mdr_data_out[113])
         ) ;
    xnor2 ix31157 (.Y (nx31156), .A0 (nx12894), .A1 (nx13298)) ;
    oai22 ix12895 (.Y (nx12894), .A0 (nx31146), .A1 (nx31159), .B0 (nx31166), .B1 (
          nx35537)) ;
    aoi32 ix31162 (.Y (nx31161), .A0 (nx12876), .A1 (nx35025), .A2 (nx31164), .B0 (
          mdr_data_out[114]), .B1 (nx35019)) ;
    oai21 ix12877 (.Y (nx12876), .A0 (mdr_data_out[112]), .A1 (mdr_data_out[113]
          ), .B0 (mdr_data_out[114])) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_18), .QB (nx31166), .D (nx22033)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22024 (.Y (nx22023), .A0 (nx31171), .A1 (nx35525), .B0 (nx31173)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_19), .QB (nx31171), .D (nx22023)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31174 (.Y (nx31173), .A0 (nx35533), .A1 (nx13326), .A2 (nx36163)) ;
    xnor2 ix13327 (.Y (nx13326), .A0 (nx31176), .A1 (nx13299)) ;
    aoi22 ix31177 (.Y (nx31176), .A0 (booth_booth_integrtaion_6_booth_output_19)
          , .A1 (nx12914), .B0 (nx12894), .B1 (nx13298)) ;
    nor02ii ix31180 (.Y (nx31179), .A0 (nx12880), .A1 (mdr_data_out[115])) ;
    nor03_2x ix12881 (.Y (nx12880), .A0 (mdr_data_out[114]), .A1 (
             mdr_data_out[112]), .A2 (mdr_data_out[113])) ;
    nor04 ix12905 (.Y (nx12904), .A0 (mdr_data_out[115]), .A1 (mdr_data_out[114]
          ), .A2 (mdr_data_out[112]), .A3 (mdr_data_out[113])) ;
    xnor2 ix31194 (.Y (nx31193), .A0 (nx12942), .A1 (nx13300)) ;
    oai22 ix12943 (.Y (nx12942), .A0 (nx31176), .A1 (nx31196), .B0 (nx31205), .B1 (
          nx35539)) ;
    aoi32 ix31199 (.Y (nx31198), .A0 (nx12924), .A1 (nx35025), .A2 (nx31203), .B0 (
          mdr_data_out[116]), .B1 (nx35019)) ;
    nand02 ix12925 (.Y (nx12924), .A0 (nx31201), .A1 (mdr_data_out[116])) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_20), .QB (nx31205), .D (nx22013)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22004 (.Y (nx22003), .A0 (nx31210), .A1 (nx35525), .B0 (nx31212)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_21), .QB (nx31210), .D (nx22003)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31213 (.Y (nx31212), .A0 (nx35533), .A1 (nx13302), .A2 (nx36163)) ;
    xnor2 ix13303 (.Y (nx13302), .A0 (nx31215), .A1 (nx13301)) ;
    aoi22 ix31216 (.Y (nx31215), .A0 (booth_booth_integrtaion_6_booth_output_21)
          , .A1 (nx12962), .B0 (nx12942), .B1 (nx13300)) ;
    nor02ii ix31219 (.Y (nx31218), .A0 (nx12928), .A1 (mdr_data_out[117])) ;
    nor02ii ix12929 (.Y (nx12928), .A0 (mdr_data_out[116]), .A1 (nx12904)) ;
    nor02ii ix12953 (.Y (nx12952), .A0 (mdr_data_out[117]), .A1 (nx12928)) ;
    xnor2 ix31229 (.Y (nx31228), .A0 (nx12990), .A1 (nx13303)) ;
    oai22 ix12991 (.Y (nx12990), .A0 (nx31215), .A1 (nx31231), .B0 (nx31240), .B1 (
          nx35541)) ;
    aoi32 ix31234 (.Y (nx31233), .A0 (nx12972), .A1 (nx35025), .A2 (nx31238), .B0 (
          mdr_data_out[118]), .B1 (nx35019)) ;
    nand02 ix12973 (.Y (nx12972), .A0 (nx31236), .A1 (mdr_data_out[118])) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_22), .QB (nx31240), .D (nx21993)
         , .CLK (clk), .R (rst)) ;
    oai21 ix21984 (.Y (nx21983), .A0 (nx31245), .A1 (nx35525), .B0 (nx31247)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_23), .QB (nx31245), .D (nx21983)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31248 (.Y (nx31247), .A0 (nx35533), .A1 (nx13278), .A2 (nx35527)) ;
    xnor2 ix13279 (.Y (nx13278), .A0 (nx31250), .A1 (nx13305)) ;
    aoi22 ix31251 (.Y (nx31250), .A0 (booth_booth_integrtaion_6_booth_output_23)
          , .A1 (nx13010), .B0 (nx12990), .B1 (nx13303)) ;
    nor02ii ix31254 (.Y (nx31253), .A0 (nx12976), .A1 (mdr_data_out[119])) ;
    nor02ii ix12977 (.Y (nx12976), .A0 (mdr_data_out[118]), .A1 (nx12952)) ;
    nor02ii ix13001 (.Y (nx13000), .A0 (mdr_data_out[119]), .A1 (nx12976)) ;
    xnor2 ix31264 (.Y (nx31263), .A0 (nx13038), .A1 (nx13307)) ;
    oai22 ix13039 (.Y (nx13038), .A0 (nx31250), .A1 (nx31266), .B0 (nx31275), .B1 (
          nx35543)) ;
    aoi32 ix31269 (.Y (nx31268), .A0 (nx13020), .A1 (nx35025), .A2 (nx31273), .B0 (
          mdr_data_out[120]), .B1 (nx35019)) ;
    nand02 ix13021 (.Y (nx13020), .A0 (nx31271), .A1 (mdr_data_out[120])) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_24), .QB (nx31275), .D (nx21973)
         , .CLK (clk), .R (rst)) ;
    oai21 ix21964 (.Y (nx21963), .A0 (nx31280), .A1 (nx35527), .B0 (nx31282)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_25), .QB (nx31280), .D (nx21963)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31283 (.Y (nx31282), .A0 (nx35533), .A1 (nx13254), .A2 (nx35527)) ;
    xnor2 ix13255 (.Y (nx13254), .A0 (nx31285), .A1 (nx13308)) ;
    aoi22 ix31286 (.Y (nx31285), .A0 (booth_booth_integrtaion_6_booth_output_25)
          , .A1 (nx13058), .B0 (nx13038), .B1 (nx13307)) ;
    nor02ii ix31289 (.Y (nx31288), .A0 (nx13024), .A1 (mdr_data_out[121])) ;
    nor02ii ix13025 (.Y (nx13024), .A0 (mdr_data_out[120]), .A1 (nx13000)) ;
    nor02ii ix13049 (.Y (nx13048), .A0 (mdr_data_out[121]), .A1 (nx13024)) ;
    xnor2 ix31299 (.Y (nx31298), .A0 (nx13086), .A1 (nx13309)) ;
    oai22 ix13087 (.Y (nx13086), .A0 (nx31285), .A1 (nx31301), .B0 (nx31310), .B1 (
          nx35545)) ;
    aoi32 ix31304 (.Y (nx31303), .A0 (nx13068), .A1 (nx35025), .A2 (nx31308), .B0 (
          mdr_data_out[122]), .B1 (nx35019)) ;
    nand02 ix13069 (.Y (nx13068), .A0 (nx31306), .A1 (mdr_data_out[122])) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_26), .QB (nx31310), .D (nx21953)
         , .CLK (clk), .R (rst)) ;
    oai21 ix21944 (.Y (nx21943), .A0 (nx31315), .A1 (nx35527), .B0 (nx31317)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_27), .QB (nx31315), .D (nx21943)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31318 (.Y (nx31317), .A0 (nx35533), .A1 (nx13230), .A2 (nx35527)) ;
    xnor2 ix13231 (.Y (nx13230), .A0 (nx31320), .A1 (nx13310)) ;
    aoi22 ix31321 (.Y (nx31320), .A0 (booth_booth_integrtaion_6_booth_output_27)
          , .A1 (nx13106), .B0 (nx13086), .B1 (nx13309)) ;
    nor02ii ix31324 (.Y (nx31323), .A0 (nx13072), .A1 (mdr_data_out[123])) ;
    nor02ii ix13073 (.Y (nx13072), .A0 (mdr_data_out[122]), .A1 (nx13048)) ;
    nor02ii ix13097 (.Y (nx13096), .A0 (mdr_data_out[123]), .A1 (nx13072)) ;
    xnor2 ix31334 (.Y (nx31333), .A0 (nx13134), .A1 (nx13311)) ;
    oai22 ix13135 (.Y (nx13134), .A0 (nx31320), .A1 (nx31336), .B0 (nx31345), .B1 (
          nx35547)) ;
    aoi32 ix31339 (.Y (nx31338), .A0 (nx13116), .A1 (nx35025), .A2 (nx31343), .B0 (
          mdr_data_out[124]), .B1 (nx35019)) ;
    nand02 ix13117 (.Y (nx13116), .A0 (nx31341), .A1 (mdr_data_out[124])) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_28), .QB (nx31345), .D (nx21933)
         , .CLK (clk), .R (rst)) ;
    oai21 ix21924 (.Y (nx21923), .A0 (nx31350), .A1 (nx35527), .B0 (nx31352)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_29), .QB (nx31350), .D (nx21923)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31353 (.Y (nx31352), .A0 (nx36171), .A1 (nx13206), .A2 (nx35527)) ;
    xnor2 ix13207 (.Y (nx13206), .A0 (nx31355), .A1 (nx13312)) ;
    aoi22 ix31356 (.Y (nx31355), .A0 (booth_booth_integrtaion_6_booth_output_29)
          , .A1 (nx13154), .B0 (nx13134), .B1 (nx13311)) ;
    nor02ii ix31359 (.Y (nx31358), .A0 (nx13120), .A1 (mdr_data_out[125])) ;
    nor02ii ix13121 (.Y (nx13120), .A0 (mdr_data_out[124]), .A1 (nx13096)) ;
    nor02ii ix13145 (.Y (nx13144), .A0 (mdr_data_out[125]), .A1 (nx13120)) ;
    xnor2 ix31369 (.Y (nx31368), .A0 (nx13182), .A1 (nx13192)) ;
    oai22 ix13183 (.Y (nx13182), .A0 (nx31355), .A1 (nx31371), .B0 (nx31380), .B1 (
          nx35549)) ;
    aoi32 ix31374 (.Y (nx31373), .A0 (nx13164), .A1 (nx35027), .A2 (nx31378), .B0 (
          mdr_data_out[126]), .B1 (nx35021)) ;
    nand02 ix13165 (.Y (nx13164), .A0 (nx31376), .A1 (mdr_data_out[126])) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_31), .QB (nx31380), .D (nx21913)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix31384 (.Y (nx31383), .A0 (mdr_data_out[127]), .A1 (nx35021), .B0 (
          nx35027), .B1 (nx13184)) ;
    xnor2 ix13185 (.Y (nx13184), .A0 (mdr_data_out[127]), .A1 (nx13168)) ;
    nor02ii ix13169 (.Y (nx13168), .A0 (mdr_data_out[126]), .A1 (nx13144)) ;
    aoi32 ix31388 (.Y (nx31387), .A0 (nx13140), .A1 (nx35027), .A2 (nx31376), .B0 (
          mdr_data_out[125]), .B1 (nx35021)) ;
    aoi32 ix31391 (.Y (nx31390), .A0 (nx13092), .A1 (nx35027), .A2 (nx31341), .B0 (
          mdr_data_out[123]), .B1 (nx35021)) ;
    aoi32 ix31394 (.Y (nx31393), .A0 (nx13044), .A1 (nx35027), .A2 (nx31306), .B0 (
          mdr_data_out[121]), .B1 (nx35021)) ;
    aoi32 ix31397 (.Y (nx31396), .A0 (nx12996), .A1 (nx35027), .A2 (nx31271), .B0 (
          mdr_data_out[119]), .B1 (nx35021)) ;
    aoi32 ix31400 (.Y (nx31399), .A0 (nx12948), .A1 (nx35027), .A2 (nx31236), .B0 (
          mdr_data_out[117]), .B1 (nx35021)) ;
    aoi32 ix31403 (.Y (nx31402), .A0 (nx12900), .A1 (nx12836), .A2 (nx31201), .B0 (
          mdr_data_out[115]), .B1 (nx35023)) ;
    aoi32 ix31406 (.Y (nx31405), .A0 (nx12850), .A1 (nx12836), .A2 (nx31150), .B0 (
          mdr_data_out[113]), .B1 (nx35023)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_6_booth_output_16), .QB (nx31131), .D (nx22053)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_6_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_6_15), .QB (nx31409), .D (nx22063), .CLK (
         clk), .R (rst)) ;
    aoi21 ix13575 (.Y (nx13574), .A0 (label_7_output[0]), .A1 (nx35771), .B0 (
          nx35919)) ;
    oai21 ix23624 (.Y (nx23623), .A0 (nx31429), .A1 (nx34785), .B0 (nx31431)) ;
    dff max_calc_reg_comparator_fourth_inp2_0 (.Q (\$dummy [468]), .QB (nx31429)
        , .D (nx23623), .CLK (clk)) ;
    nand03 ix31432 (.Y (nx31431), .A0 (label_8_output[0]), .A1 (nx35461), .A2 (
           nx34785)) ;
    dffr labelsregfile_label8_loop1_0_fx_reg_q (.Q (label_8_output[0]), .QB (
         \$dummy [469]), .D (nx23073), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_0 (.Q (label_8_input_0), .D (nx14902), .CLK (nx34529
          )) ;
    oai21 ix14903 (.Y (nx14902), .A0 (nx31437), .A1 (nx34429), .B0 (nx31441)) ;
    dffr reg_label_8_input_state_machine_0 (.Q (label_8_input_state_machine_0), 
         .QB (nx31437), .D (nx23063), .CLK (clk), .R (rst)) ;
    oai21 ix31442 (.Y (nx31441), .A0 (nx35775), .A1 (label_8_output[0]), .B0 (
          nx14890)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integration_output_7_1), .QB (\$dummy [470]), .D (nx23043)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integration_output_7_2), .QB (nx31862), .D (nx23033), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integration_output_7_3), .QB (\$dummy [471]), .D (nx23023)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integration_output_7_4), .QB (nx31860), .D (nx23013), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integration_output_7_5), .QB (\$dummy [472]), .D (nx23003)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integration_output_7_6), .QB (nx31858), .D (nx22993), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integration_output_7_7), .QB (\$dummy [473]), .D (nx22983)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integration_output_7_8), .QB (nx31856), .D (nx22973), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_10_fx_reg_q (.Q (
         booth_booth_integration_output_7_9), .QB (\$dummy [474]), .D (nx22963)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_11_fx_reg_q (.Q (
         booth_booth_integration_output_7_10), .QB (nx31854), .D (nx22953), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_12_fx_reg_q (.Q (
         booth_booth_integration_output_7_11), .QB (\$dummy [475]), .D (nx22943)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_13_fx_reg_q (.Q (
         booth_booth_integration_output_7_12), .QB (nx31852), .D (nx22933), .CLK (
         clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_14_fx_reg_q (.Q (
         booth_booth_integration_output_7_13), .QB (\$dummy [476]), .D (nx22923)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_15_fx_reg_q (.Q (
         booth_booth_integration_output_7_14), .QB (nx31850), .D (nx22913), .CLK (
         clk), .R (rst)) ;
    aoi22 ix31491 (.Y (nx31490), .A0 (mdr_data_out[15]), .A1 (nx35043), .B0 (
          nx14688), .B1 (nx14694)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_0_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_reg_output_0), .QB (\$dummy [477]), .D (
         nx22553), .CLK (clk), .R (rst)) ;
    dffs_ni booth_booth_integrtaion_7_shift_Reg_reg_count_0 (.Q (
            booth_booth_integrtaion_7_shift_Reg_count_0), .QB (\$dummy [478]), .D (
            nx22539), .CLK (clk), .S (nx34493)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_9_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_reg_output_9), .QB (\$dummy [479]), .D (
         nx22733), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_9 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_9), .QB (\$dummy [480]), .D (
         nx22723), .CLK (clk), .R (nx34493)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_8_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_8), .QB (\$dummy [481]), .D (
         nx22713), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_8 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_8), .QB (\$dummy [482]), .D (
         nx22703), .CLK (clk), .R (nx34493)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_7_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_7), .QB (\$dummy [483]), .D (
         nx22693), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_7 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_7), .QB (\$dummy [484]), .D (
         nx22683), .CLK (clk), .R (nx34493)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_6_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_6), .QB (\$dummy [485]), .D (
         nx22673), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_6 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_6), .QB (\$dummy [486]), .D (
         nx22663), .CLK (clk), .R (nx34491)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_5_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_5), .QB (\$dummy [487]), .D (
         nx22653), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_5 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_5), .QB (\$dummy [488]), .D (
         nx22643), .CLK (clk), .R (nx34491)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_4_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_4), .QB (\$dummy [489]), .D (
         nx22633), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_4 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_4), .QB (\$dummy [490]), .D (
         nx22623), .CLK (clk), .R (nx34491)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_3_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_3), .QB (\$dummy [491]), .D (
         nx22613), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_3 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_3), .QB (\$dummy [492]), .D (
         nx22603), .CLK (clk), .R (nx34491)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_2_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_2), .QB (\$dummy [493]), .D (
         nx22593), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_2 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_2), .QB (\$dummy [494]), .D (
         nx22583), .CLK (clk), .R (nx34491)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_Reg_loop1_1_fx_reg_q (.Q (
         booth_booth_integrtaion_7_shift_Reg_output_1), .QB (\$dummy [495]), .D (
         nx22573), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_shift_Reg_reg_count_1 (.Q (
         booth_booth_integrtaion_7_shift_Reg_count_1), .QB (\$dummy [496]), .D (
         nx22563), .CLK (clk), .R (nx34491)) ;
    nand02 ix22534 (.Y (nx22533), .A0 (nx35839), .A1 (nx35029)) ;
    dffs_ni booth_booth_integrtaion_7_shift_Reg_reg_en (.Q (\$dummy [497]), .QB (
            nx31537), .D (nx22533), .CLK (clk), .S (nx34491)) ;
    nand02 ix14689 (.Y (nx14688), .A0 (nx31558), .A1 (nx31570)) ;
    oai21 ix31559 (.Y (nx31558), .A0 (nx35057), .A1 (nx35051), .B0 (
          mdr_data_out[128])) ;
    oai21 ix22744 (.Y (nx22743), .A0 (nx31563), .A1 (nx35551), .B0 (nx31565)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_0_fx_reg_q (.Q (\$dummy [498]), .QB (
         nx31563), .D (nx22743), .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_1_fx_reg_q (.Q (\$dummy [499]), .QB (
         nx31567), .D (nx23053), .CLK (clk), .R (rst)) ;
    xnor2 ix31575 (.Y (nx31574), .A0 (nx14158), .A1 (nx13334)) ;
    oai21 ix22884 (.Y (nx22883), .A0 (nx31580), .A1 (nx35551), .B0 (nx31582)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_18_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_17), .QB (nx31580), .D (nx22883)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31583 (.Y (nx31582), .A0 (nx35559), .A1 (nx14666), .A2 (nx36179)) ;
    xnor2 ix14667 (.Y (nx14666), .A0 (nx31585), .A1 (nx13335)) ;
    aoi22 ix31586 (.Y (nx31585), .A0 (booth_booth_integrtaion_7_booth_output_17)
          , .A1 (nx14182), .B0 (nx14158), .B1 (nx13334)) ;
    nand02 ix14167 (.Y (nx14166), .A0 (mdr_data_out[129]), .A1 (
           mdr_data_out[128])) ;
    or02 ix31590 (.Y (nx31589), .A0 (mdr_data_out[128]), .A1 (mdr_data_out[129])
         ) ;
    xnor2 ix31596 (.Y (nx31595), .A0 (nx14210), .A1 (nx13336)) ;
    oai22 ix14211 (.Y (nx14210), .A0 (nx31585), .A1 (nx31598), .B0 (nx31605), .B1 (
          nx35563)) ;
    aoi32 ix31601 (.Y (nx31600), .A0 (nx14192), .A1 (nx35057), .A2 (nx31603), .B0 (
          mdr_data_out[130]), .B1 (nx35051)) ;
    oai21 ix14193 (.Y (nx14192), .A0 (mdr_data_out[128]), .A1 (mdr_data_out[129]
          ), .B0 (mdr_data_out[130])) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_19_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_18), .QB (nx31605), .D (nx22873)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22864 (.Y (nx22863), .A0 (nx31610), .A1 (nx35551), .B0 (nx31612)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_20_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_19), .QB (nx31610), .D (nx22863)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31613 (.Y (nx31612), .A0 (nx35559), .A1 (nx14642), .A2 (nx36179)) ;
    xnor2 ix14643 (.Y (nx14642), .A0 (nx31615), .A1 (nx13337)) ;
    aoi22 ix31616 (.Y (nx31615), .A0 (booth_booth_integrtaion_7_booth_output_19)
          , .A1 (nx14230), .B0 (nx14210), .B1 (nx13336)) ;
    nor02ii ix31619 (.Y (nx31618), .A0 (nx14196), .A1 (mdr_data_out[131])) ;
    nor03_2x ix14197 (.Y (nx14196), .A0 (mdr_data_out[130]), .A1 (
             mdr_data_out[128]), .A2 (mdr_data_out[129])) ;
    nor04 ix14221 (.Y (nx14220), .A0 (mdr_data_out[131]), .A1 (mdr_data_out[130]
          ), .A2 (mdr_data_out[128]), .A3 (mdr_data_out[129])) ;
    xnor2 ix31633 (.Y (nx31632), .A0 (nx14258), .A1 (nx13339)) ;
    oai22 ix14259 (.Y (nx14258), .A0 (nx31615), .A1 (nx31635), .B0 (nx31644), .B1 (
          nx35565)) ;
    aoi32 ix31638 (.Y (nx31637), .A0 (nx14240), .A1 (nx35057), .A2 (nx31642), .B0 (
          mdr_data_out[132]), .B1 (nx35051)) ;
    nand02 ix14241 (.Y (nx14240), .A0 (nx31640), .A1 (mdr_data_out[132])) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_21_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_20), .QB (nx31644), .D (nx22853)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22844 (.Y (nx22843), .A0 (nx31649), .A1 (nx35551), .B0 (nx31651)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_22_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_21), .QB (nx31649), .D (nx22843)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31652 (.Y (nx31651), .A0 (nx35559), .A1 (nx14618), .A2 (nx36179)) ;
    xnor2 ix14619 (.Y (nx14618), .A0 (nx31654), .A1 (nx13341)) ;
    aoi22 ix31655 (.Y (nx31654), .A0 (booth_booth_integrtaion_7_booth_output_21)
          , .A1 (nx14278), .B0 (nx14258), .B1 (nx13339)) ;
    nor02ii ix31658 (.Y (nx31657), .A0 (nx14244), .A1 (mdr_data_out[133])) ;
    nor02ii ix14245 (.Y (nx14244), .A0 (mdr_data_out[132]), .A1 (nx14220)) ;
    nor02ii ix14269 (.Y (nx14268), .A0 (mdr_data_out[133]), .A1 (nx14244)) ;
    xnor2 ix31668 (.Y (nx31667), .A0 (nx14306), .A1 (nx13343)) ;
    oai22 ix14307 (.Y (nx14306), .A0 (nx31654), .A1 (nx31670), .B0 (nx31679), .B1 (
          nx35567)) ;
    aoi32 ix31673 (.Y (nx31672), .A0 (nx14288), .A1 (nx35057), .A2 (nx31677), .B0 (
          mdr_data_out[134]), .B1 (nx35051)) ;
    nand02 ix14289 (.Y (nx14288), .A0 (nx31675), .A1 (mdr_data_out[134])) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_23_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_22), .QB (nx31679), .D (nx22833)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22824 (.Y (nx22823), .A0 (nx31684), .A1 (nx35551), .B0 (nx31686)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_24_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_23), .QB (nx31684), .D (nx22823)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31687 (.Y (nx31686), .A0 (nx35559), .A1 (nx14594), .A2 (nx35553)) ;
    xnor2 ix14595 (.Y (nx14594), .A0 (nx31689), .A1 (nx13344)) ;
    aoi22 ix31690 (.Y (nx31689), .A0 (booth_booth_integrtaion_7_booth_output_23)
          , .A1 (nx14326), .B0 (nx14306), .B1 (nx13343)) ;
    nor02ii ix31693 (.Y (nx31692), .A0 (nx14292), .A1 (mdr_data_out[135])) ;
    nor02ii ix14293 (.Y (nx14292), .A0 (mdr_data_out[134]), .A1 (nx14268)) ;
    nor02ii ix14317 (.Y (nx14316), .A0 (mdr_data_out[135]), .A1 (nx14292)) ;
    xnor2 ix31703 (.Y (nx31702), .A0 (nx14354), .A1 (nx13345)) ;
    oai22 ix14355 (.Y (nx14354), .A0 (nx31689), .A1 (nx31705), .B0 (nx31714), .B1 (
          nx35569)) ;
    aoi32 ix31708 (.Y (nx31707), .A0 (nx14336), .A1 (nx35057), .A2 (nx31712), .B0 (
          mdr_data_out[136]), .B1 (nx35051)) ;
    nand02 ix14337 (.Y (nx14336), .A0 (nx31710), .A1 (mdr_data_out[136])) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_25_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_24), .QB (nx31714), .D (nx22813)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22804 (.Y (nx22803), .A0 (nx31719), .A1 (nx35553), .B0 (nx31721)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_26_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_25), .QB (nx31719), .D (nx22803)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31722 (.Y (nx31721), .A0 (nx35559), .A1 (nx14570), .A2 (nx35553)) ;
    xnor2 ix14571 (.Y (nx14570), .A0 (nx31724), .A1 (nx13346)) ;
    aoi22 ix31725 (.Y (nx31724), .A0 (booth_booth_integrtaion_7_booth_output_25)
          , .A1 (nx14374), .B0 (nx14354), .B1 (nx13345)) ;
    nor02ii ix31728 (.Y (nx31727), .A0 (nx14340), .A1 (mdr_data_out[137])) ;
    nor02ii ix14341 (.Y (nx14340), .A0 (mdr_data_out[136]), .A1 (nx14316)) ;
    nor02ii ix14365 (.Y (nx14364), .A0 (mdr_data_out[137]), .A1 (nx14340)) ;
    xnor2 ix31738 (.Y (nx31737), .A0 (nx14402), .A1 (nx13347)) ;
    oai22 ix14403 (.Y (nx14402), .A0 (nx31724), .A1 (nx31740), .B0 (nx31749), .B1 (
          nx35571)) ;
    aoi32 ix31743 (.Y (nx31742), .A0 (nx14384), .A1 (nx35057), .A2 (nx31747), .B0 (
          mdr_data_out[138]), .B1 (nx35051)) ;
    nand02 ix14385 (.Y (nx14384), .A0 (nx31745), .A1 (mdr_data_out[138])) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_27_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_26), .QB (nx31749), .D (nx22793)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22784 (.Y (nx22783), .A0 (nx31754), .A1 (nx35553), .B0 (nx31756)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_28_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_27), .QB (nx31754), .D (nx22783)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31757 (.Y (nx31756), .A0 (nx35559), .A1 (nx14546), .A2 (nx35553)) ;
    xnor2 ix14547 (.Y (nx14546), .A0 (nx31759), .A1 (nx13348)) ;
    aoi22 ix31760 (.Y (nx31759), .A0 (booth_booth_integrtaion_7_booth_output_27)
          , .A1 (nx14422), .B0 (nx14402), .B1 (nx13347)) ;
    nor02ii ix31763 (.Y (nx31762), .A0 (nx14388), .A1 (mdr_data_out[139])) ;
    nor02ii ix14389 (.Y (nx14388), .A0 (mdr_data_out[138]), .A1 (nx14364)) ;
    nor02ii ix14413 (.Y (nx14412), .A0 (mdr_data_out[139]), .A1 (nx14388)) ;
    xnor2 ix31773 (.Y (nx31772), .A0 (nx14450), .A1 (nx13349)) ;
    oai22 ix14451 (.Y (nx14450), .A0 (nx31759), .A1 (nx31775), .B0 (nx31784), .B1 (
          nx35573)) ;
    aoi32 ix31778 (.Y (nx31777), .A0 (nx14432), .A1 (nx35057), .A2 (nx31782), .B0 (
          mdr_data_out[140]), .B1 (nx35051)) ;
    nand02 ix14433 (.Y (nx14432), .A0 (nx31780), .A1 (mdr_data_out[140])) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_29_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_28), .QB (nx31784), .D (nx22773)
         , .CLK (clk), .R (rst)) ;
    oai21 ix22764 (.Y (nx22763), .A0 (nx31789), .A1 (nx35553), .B0 (nx31791)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_30_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_29), .QB (nx31789), .D (nx22763)
         , .CLK (clk), .R (rst)) ;
    nand03 ix31792 (.Y (nx31791), .A0 (nx36187), .A1 (nx14522), .A2 (nx35553)) ;
    xnor2 ix14523 (.Y (nx14522), .A0 (nx31794), .A1 (nx13351)) ;
    aoi22 ix31795 (.Y (nx31794), .A0 (booth_booth_integrtaion_7_booth_output_29)
          , .A1 (nx14470), .B0 (nx14450), .B1 (nx13349)) ;
    nor02ii ix31798 (.Y (nx31797), .A0 (nx14436), .A1 (mdr_data_out[141])) ;
    nor02ii ix14437 (.Y (nx14436), .A0 (mdr_data_out[140]), .A1 (nx14412)) ;
    nor02ii ix14461 (.Y (nx14460), .A0 (mdr_data_out[141]), .A1 (nx14436)) ;
    xnor2 ix31808 (.Y (nx31807), .A0 (nx14498), .A1 (nx14508)) ;
    oai22 ix14499 (.Y (nx14498), .A0 (nx31794), .A1 (nx31810), .B0 (nx31819), .B1 (
          nx35575)) ;
    aoi32 ix31813 (.Y (nx31812), .A0 (nx14480), .A1 (nx35059), .A2 (nx31817), .B0 (
          mdr_data_out[142]), .B1 (nx35053)) ;
    nand02 ix14481 (.Y (nx14480), .A0 (nx31815), .A1 (mdr_data_out[142])) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_32_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_31), .QB (nx31819), .D (nx22753)
         , .CLK (clk), .R (rst)) ;
    aoi22 ix31823 (.Y (nx31822), .A0 (mdr_data_out[143]), .A1 (nx35053), .B0 (
          nx35059), .B1 (nx14500)) ;
    xnor2 ix14501 (.Y (nx14500), .A0 (mdr_data_out[143]), .A1 (nx14484)) ;
    nor02ii ix14485 (.Y (nx14484), .A0 (mdr_data_out[142]), .A1 (nx14460)) ;
    aoi32 ix31827 (.Y (nx31826), .A0 (nx14456), .A1 (nx35059), .A2 (nx31815), .B0 (
          mdr_data_out[141]), .B1 (nx35053)) ;
    aoi32 ix31830 (.Y (nx31829), .A0 (nx14408), .A1 (nx35059), .A2 (nx31780), .B0 (
          mdr_data_out[139]), .B1 (nx35053)) ;
    aoi32 ix31833 (.Y (nx31832), .A0 (nx14360), .A1 (nx35059), .A2 (nx31745), .B0 (
          mdr_data_out[137]), .B1 (nx35053)) ;
    aoi32 ix31836 (.Y (nx31835), .A0 (nx14312), .A1 (nx35059), .A2 (nx31710), .B0 (
          mdr_data_out[135]), .B1 (nx35053)) ;
    aoi32 ix31839 (.Y (nx31838), .A0 (nx14264), .A1 (nx35059), .A2 (nx31675), .B0 (
          mdr_data_out[133]), .B1 (nx35053)) ;
    aoi32 ix31842 (.Y (nx31841), .A0 (nx14216), .A1 (nx14152), .A2 (nx31640), .B0 (
          mdr_data_out[131]), .B1 (nx35055)) ;
    aoi32 ix31845 (.Y (nx31844), .A0 (nx14166), .A1 (nx14152), .A2 (nx31589), .B0 (
          mdr_data_out[129]), .B1 (nx35055)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_17_fx_reg_q (.Q (
         booth_booth_integrtaion_7_booth_output_16), .QB (nx31570), .D (nx22893)
         , .CLK (clk), .R (rst)) ;
    dffr booth_booth_integrtaion_7_p_Reg_loop1_16_fx_reg_q (.Q (
         booth_booth_integration_output_7_15), .QB (nx31848), .D (nx22903), .CLK (
         clk), .R (rst)) ;
    aoi21 ix14891 (.Y (nx14890), .A0 (label_8_output[0]), .A1 (nx35775), .B0 (
          nx35919)) ;
    xnor2 ix15875 (.Y (nx15874), .A0 (nx31867), .A1 (nx15872)) ;
    aoi22 ix31868 (.Y (nx31867), .A0 (nx31869), .A1 (
          max_calc_comparator_fourth_inp1_14), .B0 (nx15360), .B1 (nx15778)) ;
    dff max_calc_reg_comparator_fourth_inp2_14 (.Q (\$dummy [500]), .QB (nx31869
        ), .D (nx23353), .CLK (clk)) ;
    oai21 ix23354 (.Y (nx23353), .A0 (nx31869), .A1 (nx34785), .B0 (nx31872)) ;
    dffr labelsregfile_label8_loop1_14_fx_reg_q (.Q (label_8_output[14]), .QB (
         nx32056), .D (nx23343), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_14 (.Q (label_8_input_14), .D (nx15338), .CLK (
          nx34533)) ;
    dffr reg_label_8_input_state_machine_14 (.Q (label_8_input_state_machine_14)
         , .QB (\$dummy [501]), .D (nx22523), .CLK (clk), .R (rst)) ;
    xor2 ix15335 (.Y (nx15334), .A0 (nx31882), .A1 (nx32054)) ;
    aoi22 ix31883 (.Y (nx31882), .A0 (label_8_output[13]), .A1 (
          booth_booth_integration_output_7_13), .B0 (nx15298), .B1 (nx13370)) ;
    dffr labelsregfile_label8_loop1_13_fx_reg_q (.Q (label_8_output[13]), .QB (
         \$dummy [502]), .D (nx23333), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_13 (.Q (label_8_input_13), .D (nx15312), .CLK (
          nx34533)) ;
    dffr reg_label_8_input_state_machine_13 (.Q (label_8_input_state_machine_13)
         , .QB (\$dummy [503]), .D (nx23323), .CLK (clk), .R (rst)) ;
    xnor2 ix15309 (.Y (nx15308), .A0 (nx15298), .A1 (nx32050)) ;
    oai22 ix15299 (.Y (nx15298), .A0 (nx31893), .A1 (nx32039), .B0 (nx32049), .B1 (
          nx31852)) ;
    aoi22 ix31894 (.Y (nx31893), .A0 (label_8_output[11]), .A1 (
          booth_booth_integration_output_7_11), .B0 (nx15234), .B1 (nx13368)) ;
    dffr labelsregfile_label8_loop1_11_fx_reg_q (.Q (label_8_output[11]), .QB (
         \$dummy [504]), .D (nx23293), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_11 (.Q (label_8_input_11), .D (nx15248), .CLK (
          nx34533)) ;
    dffr reg_label_8_input_state_machine_11 (.Q (label_8_input_state_machine_11)
         , .QB (\$dummy [505]), .D (nx23283), .CLK (clk), .R (rst)) ;
    xnor2 ix15245 (.Y (nx15244), .A0 (nx15234), .A1 (nx32035)) ;
    oai22 ix15235 (.Y (nx15234), .A0 (nx31904), .A1 (nx32024), .B0 (nx32034), .B1 (
          nx31854)) ;
    aoi22 ix31905 (.Y (nx31904), .A0 (label_8_output[9]), .A1 (
          booth_booth_integration_output_7_9), .B0 (nx15170), .B1 (nx13365)) ;
    dffr labelsregfile_label8_loop1_9_fx_reg_q (.Q (label_8_output[9]), .QB (
         \$dummy [506]), .D (nx23253), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_9 (.Q (label_8_input_9), .D (nx15184), .CLK (nx34533
          )) ;
    dffr reg_label_8_input_state_machine_9 (.Q (label_8_input_state_machine_9), 
         .QB (\$dummy [507]), .D (nx23243), .CLK (clk), .R (rst)) ;
    xnor2 ix15181 (.Y (nx15180), .A0 (nx15170), .A1 (nx32020)) ;
    oai22 ix15171 (.Y (nx15170), .A0 (nx31915), .A1 (nx32009), .B0 (nx32019), .B1 (
          nx31856)) ;
    aoi22 ix31916 (.Y (nx31915), .A0 (label_8_output[7]), .A1 (
          booth_booth_integration_output_7_7), .B0 (nx15106), .B1 (nx13361)) ;
    dffr labelsregfile_label8_loop1_7_fx_reg_q (.Q (label_8_output[7]), .QB (
         \$dummy [508]), .D (nx23213), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_7 (.Q (label_8_input_7), .D (nx15120), .CLK (nx34531
          )) ;
    dffr reg_label_8_input_state_machine_7 (.Q (label_8_input_state_machine_7), 
         .QB (\$dummy [509]), .D (nx23203), .CLK (clk), .R (rst)) ;
    xnor2 ix15117 (.Y (nx15116), .A0 (nx15106), .A1 (nx32005)) ;
    oai22 ix15107 (.Y (nx15106), .A0 (nx31926), .A1 (nx31994), .B0 (nx32004), .B1 (
          nx31858)) ;
    aoi22 ix31927 (.Y (nx31926), .A0 (label_8_output[5]), .A1 (
          booth_booth_integration_output_7_5), .B0 (nx15042), .B1 (nx13359)) ;
    dffr labelsregfile_label8_loop1_5_fx_reg_q (.Q (label_8_output[5]), .QB (
         \$dummy [510]), .D (nx23173), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_5 (.Q (label_8_input_5), .D (nx15056), .CLK (nx34531
          )) ;
    dffr reg_label_8_input_state_machine_5 (.Q (label_8_input_state_machine_5), 
         .QB (\$dummy [511]), .D (nx23163), .CLK (clk), .R (rst)) ;
    xnor2 ix15053 (.Y (nx15052), .A0 (nx15042), .A1 (nx31990)) ;
    oai22 ix15043 (.Y (nx15042), .A0 (nx31937), .A1 (nx31979), .B0 (nx31989), .B1 (
          nx31860)) ;
    aoi22 ix31938 (.Y (nx31937), .A0 (label_8_output[3]), .A1 (
          booth_booth_integration_output_7_3), .B0 (nx14978), .B1 (nx13357)) ;
    dffr labelsregfile_label8_loop1_3_fx_reg_q (.Q (label_8_output[3]), .QB (
         \$dummy [512]), .D (nx23133), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_3 (.Q (label_8_input_3), .D (nx14992), .CLK (nx34531
          )) ;
    dffr reg_label_8_input_state_machine_3 (.Q (label_8_input_state_machine_3), 
         .QB (\$dummy [513]), .D (nx23123), .CLK (clk), .R (rst)) ;
    xnor2 ix14989 (.Y (nx14988), .A0 (nx14978), .A1 (nx31975)) ;
    oai22 ix14979 (.Y (nx14978), .A0 (nx31948), .A1 (nx31964), .B0 (nx31974), .B1 (
          nx31862)) ;
    aoi32 ix31949 (.Y (nx31948), .A0 (label_8_output[0]), .A1 (nx35775), .A2 (
          nx13355), .B0 (label_8_output[1]), .B1 (
          booth_booth_integration_output_7_1)) ;
    dffr labelsregfile_label8_loop1_1_fx_reg_q (.Q (label_8_output[1]), .QB (
         \$dummy [514]), .D (nx23093), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_1 (.Q (label_8_input_1), .D (nx14928), .CLK (nx34531
          )) ;
    dffr reg_label_8_input_state_machine_1 (.Q (label_8_input_state_machine_1), 
         .QB (\$dummy [515]), .D (nx23083), .CLK (clk), .R (rst)) ;
    xor2 ix14925 (.Y (nx14924), .A0 (nx31959), .A1 (nx31961)) ;
    nand02 ix31960 (.Y (nx31959), .A0 (label_8_output[0]), .A1 (nx35775)) ;
    xnor2 ix31962 (.Y (nx31961), .A0 (booth_booth_integration_output_7_1), .A1 (
          label_8_output[1])) ;
    dffr labelsregfile_label8_loop1_2_fx_reg_q (.Q (label_8_output[2]), .QB (
         nx31974), .D (nx23113), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_2 (.Q (label_8_input_2), .D (nx14960), .CLK (nx34531
          )) ;
    dffr reg_label_8_input_state_machine_2 (.Q (label_8_input_state_machine_2), 
         .QB (\$dummy [516]), .D (nx23103), .CLK (clk), .R (rst)) ;
    xor2 ix14957 (.Y (nx14956), .A0 (nx31948), .A1 (nx31964)) ;
    xnor2 ix31976 (.Y (nx31975), .A0 (booth_booth_integration_output_7_3), .A1 (
          label_8_output[3])) ;
    dffr labelsregfile_label8_loop1_4_fx_reg_q (.Q (label_8_output[4]), .QB (
         nx31989), .D (nx23153), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_4 (.Q (label_8_input_4), .D (nx15024), .CLK (nx34531
          )) ;
    dffr reg_label_8_input_state_machine_4 (.Q (label_8_input_state_machine_4), 
         .QB (\$dummy [517]), .D (nx23143), .CLK (clk), .R (rst)) ;
    xor2 ix15021 (.Y (nx15020), .A0 (nx31937), .A1 (nx31979)) ;
    xnor2 ix31991 (.Y (nx31990), .A0 (booth_booth_integration_output_7_5), .A1 (
          label_8_output[5])) ;
    dffr labelsregfile_label8_loop1_6_fx_reg_q (.Q (label_8_output[6]), .QB (
         nx32004), .D (nx23193), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_6 (.Q (label_8_input_6), .D (nx15088), .CLK (nx34531
          )) ;
    dffr reg_label_8_input_state_machine_6 (.Q (label_8_input_state_machine_6), 
         .QB (\$dummy [518]), .D (nx23183), .CLK (clk), .R (rst)) ;
    xor2 ix15085 (.Y (nx15084), .A0 (nx31926), .A1 (nx31994)) ;
    xnor2 ix32006 (.Y (nx32005), .A0 (booth_booth_integration_output_7_7), .A1 (
          label_8_output[7])) ;
    dffr labelsregfile_label8_loop1_8_fx_reg_q (.Q (label_8_output[8]), .QB (
         nx32019), .D (nx23233), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_8 (.Q (label_8_input_8), .D (nx15152), .CLK (nx34533
          )) ;
    dffr reg_label_8_input_state_machine_8 (.Q (label_8_input_state_machine_8), 
         .QB (\$dummy [519]), .D (nx23223), .CLK (clk), .R (rst)) ;
    xor2 ix15149 (.Y (nx15148), .A0 (nx31915), .A1 (nx32009)) ;
    xnor2 ix32021 (.Y (nx32020), .A0 (booth_booth_integration_output_7_9), .A1 (
          label_8_output[9])) ;
    dffr labelsregfile_label8_loop1_10_fx_reg_q (.Q (label_8_output[10]), .QB (
         nx32034), .D (nx23273), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_10 (.Q (label_8_input_10), .D (nx15216), .CLK (
          nx34533)) ;
    dffr reg_label_8_input_state_machine_10 (.Q (label_8_input_state_machine_10)
         , .QB (\$dummy [520]), .D (nx23263), .CLK (clk), .R (rst)) ;
    xor2 ix15213 (.Y (nx15212), .A0 (nx31904), .A1 (nx32024)) ;
    xnor2 ix32036 (.Y (nx32035), .A0 (booth_booth_integration_output_7_11), .A1 (
          label_8_output[11])) ;
    dffr labelsregfile_label8_loop1_12_fx_reg_q (.Q (label_8_output[12]), .QB (
         nx32049), .D (nx23313), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_12 (.Q (label_8_input_12), .D (nx15280), .CLK (
          nx34533)) ;
    dffr reg_label_8_input_state_machine_12 (.Q (label_8_input_state_machine_12)
         , .QB (\$dummy [521]), .D (nx23303), .CLK (clk), .R (rst)) ;
    xor2 ix15277 (.Y (nx15276), .A0 (nx31893), .A1 (nx32039)) ;
    xnor2 ix32051 (.Y (nx32050), .A0 (booth_booth_integration_output_7_13), .A1 (
          label_8_output[13])) ;
    oai21 ix22514 (.Y (nx22513), .A0 (nx32059), .A1 (nx34785), .B0 (nx32061)) ;
    dff max_calc_reg_comparator_fourth_inp1_14 (.Q (
        max_calc_comparator_fourth_inp1_14), .QB (nx32059), .D (nx22513), .CLK (
        clk)) ;
    dffr labelsregfile_label7_loop1_14_fx_reg_q (.Q (label_7_output[14]), .QB (
         nx32245), .D (nx22503), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_14 (.Q (label_7_input_14), .D (nx14022), .CLK (
          nx34537)) ;
    dffr reg_label_7_input_state_machine_14 (.Q (label_7_input_state_machine_14)
         , .QB (\$dummy [522]), .D (nx21683), .CLK (clk), .R (rst)) ;
    xor2 ix14019 (.Y (nx14018), .A0 (nx32071), .A1 (nx32243)) ;
    aoi22 ix32072 (.Y (nx32071), .A0 (label_7_output[13]), .A1 (
          booth_booth_integration_output_6_13), .B0 (nx13982), .B1 (nx13332)) ;
    dffr labelsregfile_label7_loop1_13_fx_reg_q (.Q (label_7_output[13]), .QB (
         \$dummy [523]), .D (nx22493), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_13 (.Q (label_7_input_13), .D (nx13996), .CLK (
          nx34537)) ;
    dffr reg_label_7_input_state_machine_13 (.Q (label_7_input_state_machine_13)
         , .QB (\$dummy [524]), .D (nx22483), .CLK (clk), .R (rst)) ;
    xnor2 ix13993 (.Y (nx13992), .A0 (nx13982), .A1 (nx32239)) ;
    oai22 ix13983 (.Y (nx13982), .A0 (nx32082), .A1 (nx32228), .B0 (nx32238), .B1 (
          nx31413)) ;
    aoi22 ix32083 (.Y (nx32082), .A0 (label_7_output[11]), .A1 (
          booth_booth_integration_output_6_11), .B0 (nx13918), .B1 (nx13329)) ;
    dffr labelsregfile_label7_loop1_11_fx_reg_q (.Q (label_7_output[11]), .QB (
         \$dummy [525]), .D (nx22453), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_11 (.Q (label_7_input_11), .D (nx13932), .CLK (
          nx34537)) ;
    dffr reg_label_7_input_state_machine_11 (.Q (label_7_input_state_machine_11)
         , .QB (\$dummy [526]), .D (nx22443), .CLK (clk), .R (rst)) ;
    xnor2 ix13929 (.Y (nx13928), .A0 (nx13918), .A1 (nx32224)) ;
    oai22 ix13919 (.Y (nx13918), .A0 (nx32093), .A1 (nx32213), .B0 (nx32223), .B1 (
          nx31415)) ;
    aoi22 ix32094 (.Y (nx32093), .A0 (label_7_output[9]), .A1 (
          booth_booth_integration_output_6_9), .B0 (nx13854), .B1 (nx13325)) ;
    dffr labelsregfile_label7_loop1_9_fx_reg_q (.Q (label_7_output[9]), .QB (
         \$dummy [527]), .D (nx22413), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_9 (.Q (label_7_input_9), .D (nx13868), .CLK (nx34537
          )) ;
    dffr reg_label_7_input_state_machine_9 (.Q (label_7_input_state_machine_9), 
         .QB (\$dummy [528]), .D (nx22403), .CLK (clk), .R (rst)) ;
    xnor2 ix13865 (.Y (nx13864), .A0 (nx13854), .A1 (nx32209)) ;
    oai22 ix13855 (.Y (nx13854), .A0 (nx32104), .A1 (nx32198), .B0 (nx32208), .B1 (
          nx31417)) ;
    aoi22 ix32105 (.Y (nx32104), .A0 (label_7_output[7]), .A1 (
          booth_booth_integration_output_6_7), .B0 (nx13790), .B1 (nx13323)) ;
    dffr labelsregfile_label7_loop1_7_fx_reg_q (.Q (label_7_output[7]), .QB (
         \$dummy [529]), .D (nx22373), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_7 (.Q (label_7_input_7), .D (nx13804), .CLK (nx34535
          )) ;
    dffr reg_label_7_input_state_machine_7 (.Q (label_7_input_state_machine_7), 
         .QB (\$dummy [530]), .D (nx22363), .CLK (clk), .R (rst)) ;
    xnor2 ix13801 (.Y (nx13800), .A0 (nx13790), .A1 (nx32194)) ;
    oai22 ix13791 (.Y (nx13790), .A0 (nx32115), .A1 (nx32183), .B0 (nx32193), .B1 (
          nx31419)) ;
    aoi22 ix32116 (.Y (nx32115), .A0 (label_7_output[5]), .A1 (
          booth_booth_integration_output_6_5), .B0 (nx13726), .B1 (nx13321)) ;
    dffr labelsregfile_label7_loop1_5_fx_reg_q (.Q (label_7_output[5]), .QB (
         \$dummy [531]), .D (nx22333), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_5 (.Q (label_7_input_5), .D (nx13740), .CLK (nx34535
          )) ;
    dffr reg_label_7_input_state_machine_5 (.Q (label_7_input_state_machine_5), 
         .QB (\$dummy [532]), .D (nx22323), .CLK (clk), .R (rst)) ;
    xnor2 ix13737 (.Y (nx13736), .A0 (nx13726), .A1 (nx32179)) ;
    oai22 ix13727 (.Y (nx13726), .A0 (nx32126), .A1 (nx32168), .B0 (nx32178), .B1 (
          nx31421)) ;
    aoi22 ix32127 (.Y (nx32126), .A0 (label_7_output[3]), .A1 (
          booth_booth_integration_output_6_3), .B0 (nx13662), .B1 (nx13319)) ;
    dffr labelsregfile_label7_loop1_3_fx_reg_q (.Q (label_7_output[3]), .QB (
         \$dummy [533]), .D (nx22293), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_3 (.Q (label_7_input_3), .D (nx13676), .CLK (nx34535
          )) ;
    dffr reg_label_7_input_state_machine_3 (.Q (label_7_input_state_machine_3), 
         .QB (\$dummy [534]), .D (nx22283), .CLK (clk), .R (rst)) ;
    xnor2 ix13673 (.Y (nx13672), .A0 (nx13662), .A1 (nx32164)) ;
    oai22 ix13663 (.Y (nx13662), .A0 (nx32137), .A1 (nx32153), .B0 (nx32163), .B1 (
          nx31423)) ;
    aoi32 ix32138 (.Y (nx32137), .A0 (label_7_output[0]), .A1 (nx35771), .A2 (
          nx13315), .B0 (label_7_output[1]), .B1 (
          booth_booth_integration_output_6_1)) ;
    dffr labelsregfile_label7_loop1_1_fx_reg_q (.Q (label_7_output[1]), .QB (
         \$dummy [535]), .D (nx22253), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_1 (.Q (label_7_input_1), .D (nx13612), .CLK (nx34535
          )) ;
    dffr reg_label_7_input_state_machine_1 (.Q (label_7_input_state_machine_1), 
         .QB (\$dummy [536]), .D (nx22243), .CLK (clk), .R (rst)) ;
    xor2 ix13609 (.Y (nx13608), .A0 (nx32148), .A1 (nx32150)) ;
    nand02 ix32149 (.Y (nx32148), .A0 (label_7_output[0]), .A1 (nx35771)) ;
    xnor2 ix32151 (.Y (nx32150), .A0 (booth_booth_integration_output_6_1), .A1 (
          label_7_output[1])) ;
    dffr labelsregfile_label7_loop1_2_fx_reg_q (.Q (label_7_output[2]), .QB (
         nx32163), .D (nx22273), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_2 (.Q (label_7_input_2), .D (nx13644), .CLK (nx34535
          )) ;
    dffr reg_label_7_input_state_machine_2 (.Q (label_7_input_state_machine_2), 
         .QB (\$dummy [537]), .D (nx22263), .CLK (clk), .R (rst)) ;
    xor2 ix13641 (.Y (nx13640), .A0 (nx32137), .A1 (nx32153)) ;
    xnor2 ix32165 (.Y (nx32164), .A0 (booth_booth_integration_output_6_3), .A1 (
          label_7_output[3])) ;
    dffr labelsregfile_label7_loop1_4_fx_reg_q (.Q (label_7_output[4]), .QB (
         nx32178), .D (nx22313), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_4 (.Q (label_7_input_4), .D (nx13708), .CLK (nx34535
          )) ;
    dffr reg_label_7_input_state_machine_4 (.Q (label_7_input_state_machine_4), 
         .QB (\$dummy [538]), .D (nx22303), .CLK (clk), .R (rst)) ;
    xor2 ix13705 (.Y (nx13704), .A0 (nx32126), .A1 (nx32168)) ;
    xnor2 ix32180 (.Y (nx32179), .A0 (booth_booth_integration_output_6_5), .A1 (
          label_7_output[5])) ;
    dffr labelsregfile_label7_loop1_6_fx_reg_q (.Q (label_7_output[6]), .QB (
         nx32193), .D (nx22353), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_6 (.Q (label_7_input_6), .D (nx13772), .CLK (nx34535
          )) ;
    dffr reg_label_7_input_state_machine_6 (.Q (label_7_input_state_machine_6), 
         .QB (\$dummy [539]), .D (nx22343), .CLK (clk), .R (rst)) ;
    xor2 ix13769 (.Y (nx13768), .A0 (nx32115), .A1 (nx32183)) ;
    xnor2 ix32195 (.Y (nx32194), .A0 (booth_booth_integration_output_6_7), .A1 (
          label_7_output[7])) ;
    dffr labelsregfile_label7_loop1_8_fx_reg_q (.Q (label_7_output[8]), .QB (
         nx32208), .D (nx22393), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_8 (.Q (label_7_input_8), .D (nx13836), .CLK (nx34537
          )) ;
    dffr reg_label_7_input_state_machine_8 (.Q (label_7_input_state_machine_8), 
         .QB (\$dummy [540]), .D (nx22383), .CLK (clk), .R (rst)) ;
    xor2 ix13833 (.Y (nx13832), .A0 (nx32104), .A1 (nx32198)) ;
    xnor2 ix32210 (.Y (nx32209), .A0 (booth_booth_integration_output_6_9), .A1 (
          label_7_output[9])) ;
    dffr labelsregfile_label7_loop1_10_fx_reg_q (.Q (label_7_output[10]), .QB (
         nx32223), .D (nx22433), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_10 (.Q (label_7_input_10), .D (nx13900), .CLK (
          nx34537)) ;
    dffr reg_label_7_input_state_machine_10 (.Q (label_7_input_state_machine_10)
         , .QB (\$dummy [541]), .D (nx22423), .CLK (clk), .R (rst)) ;
    xor2 ix13897 (.Y (nx13896), .A0 (nx32093), .A1 (nx32213)) ;
    xnor2 ix32225 (.Y (nx32224), .A0 (booth_booth_integration_output_6_11), .A1 (
          label_7_output[11])) ;
    dffr labelsregfile_label7_loop1_12_fx_reg_q (.Q (label_7_output[12]), .QB (
         nx32238), .D (nx22473), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_12 (.Q (label_7_input_12), .D (nx13964), .CLK (
          nx34537)) ;
    dffr reg_label_7_input_state_machine_12 (.Q (label_7_input_state_machine_12)
         , .QB (\$dummy [542]), .D (nx22463), .CLK (clk), .R (rst)) ;
    xor2 ix13961 (.Y (nx13960), .A0 (nx32082), .A1 (nx32228)) ;
    xnor2 ix32240 (.Y (nx32239), .A0 (booth_booth_integration_output_6_13), .A1 (
          label_7_output[13])) ;
    oai22 ix15779 (.Y (nx15778), .A0 (nx32248), .A1 (nx32261), .B0 (
          max_calc_comparator_fourth_inp2_13), .B1 (nx32256)) ;
    oai21 ix23364 (.Y (nx23363), .A0 (nx32252), .A1 (nx34785), .B0 (nx32254)) ;
    dff max_calc_reg_comparator_fourth_inp2_13 (.Q (
        max_calc_comparator_fourth_inp2_13), .QB (nx32252), .D (nx23363), .CLK (
        clk)) ;
    nand03 ix32255 (.Y (nx32254), .A0 (label_8_output[13]), .A1 (nx35463), .A2 (
           nx34787)) ;
    dff max_calc_reg_comparator_fourth_inp1_13 (.Q (
        max_calc_comparator_fourth_inp1_13), .QB (nx32256), .D (nx23373), .CLK (
        clk)) ;
    oai21 ix23374 (.Y (nx23373), .A0 (nx32256), .A1 (nx34787), .B0 (nx32259)) ;
    nand03 ix32260 (.Y (nx32259), .A0 (label_7_output[13]), .A1 (nx35463), .A2 (
           nx34787)) ;
    aoi22 ix32262 (.Y (nx32261), .A0 (nx32263), .A1 (
          max_calc_comparator_fourth_inp1_12), .B0 (nx15404), .B1 (nx15762)) ;
    dff max_calc_reg_comparator_fourth_inp2_12 (.Q (\$dummy [543]), .QB (nx32263
        ), .D (nx23383), .CLK (clk)) ;
    oai21 ix23384 (.Y (nx23383), .A0 (nx32263), .A1 (nx34787), .B0 (nx32266)) ;
    oai21 ix23394 (.Y (nx23393), .A0 (nx32270), .A1 (nx34787), .B0 (nx32272)) ;
    dff max_calc_reg_comparator_fourth_inp1_12 (.Q (
        max_calc_comparator_fourth_inp1_12), .QB (nx32270), .D (nx23393), .CLK (
        clk)) ;
    oai22 ix15763 (.Y (nx15762), .A0 (nx32276), .A1 (nx32289), .B0 (
          max_calc_comparator_fourth_inp2_11), .B1 (nx32284)) ;
    oai21 ix23404 (.Y (nx23403), .A0 (nx32280), .A1 (nx34789), .B0 (nx32282)) ;
    dff max_calc_reg_comparator_fourth_inp2_11 (.Q (
        max_calc_comparator_fourth_inp2_11), .QB (nx32280), .D (nx23403), .CLK (
        clk)) ;
    nand03 ix32283 (.Y (nx32282), .A0 (label_8_output[11]), .A1 (nx35463), .A2 (
           nx34789)) ;
    dff max_calc_reg_comparator_fourth_inp1_11 (.Q (
        max_calc_comparator_fourth_inp1_11), .QB (nx32284), .D (nx23413), .CLK (
        clk)) ;
    oai21 ix23414 (.Y (nx23413), .A0 (nx32284), .A1 (nx34789), .B0 (nx32287)) ;
    nand03 ix32288 (.Y (nx32287), .A0 (label_7_output[11]), .A1 (nx35463), .A2 (
           nx34789)) ;
    aoi22 ix32290 (.Y (nx32289), .A0 (nx32291), .A1 (
          max_calc_comparator_fourth_inp1_10), .B0 (nx15448), .B1 (nx15746)) ;
    dff max_calc_reg_comparator_fourth_inp2_10 (.Q (\$dummy [544]), .QB (nx32291
        ), .D (nx23423), .CLK (clk)) ;
    oai21 ix23424 (.Y (nx23423), .A0 (nx32291), .A1 (nx34789), .B0 (nx32294)) ;
    oai21 ix23434 (.Y (nx23433), .A0 (nx32298), .A1 (nx34789), .B0 (nx32300)) ;
    dff max_calc_reg_comparator_fourth_inp1_10 (.Q (
        max_calc_comparator_fourth_inp1_10), .QB (nx32298), .D (nx23433), .CLK (
        clk)) ;
    oai22 ix15747 (.Y (nx15746), .A0 (nx32304), .A1 (nx32317), .B0 (
          max_calc_comparator_fourth_inp2_9), .B1 (nx32312)) ;
    oai21 ix23444 (.Y (nx23443), .A0 (nx32308), .A1 (nx34791), .B0 (nx32310)) ;
    dff max_calc_reg_comparator_fourth_inp2_9 (.Q (
        max_calc_comparator_fourth_inp2_9), .QB (nx32308), .D (nx23443), .CLK (
        clk)) ;
    nand03 ix32311 (.Y (nx32310), .A0 (label_8_output[9]), .A1 (nx35465), .A2 (
           nx34791)) ;
    dff max_calc_reg_comparator_fourth_inp1_9 (.Q (
        max_calc_comparator_fourth_inp1_9), .QB (nx32312), .D (nx23453), .CLK (
        clk)) ;
    oai21 ix23454 (.Y (nx23453), .A0 (nx32312), .A1 (nx34791), .B0 (nx32315)) ;
    nand03 ix32316 (.Y (nx32315), .A0 (label_7_output[9]), .A1 (nx35465), .A2 (
           nx34791)) ;
    aoi22 ix32318 (.Y (nx32317), .A0 (nx32319), .A1 (
          max_calc_comparator_fourth_inp1_8), .B0 (nx15492), .B1 (nx15730)) ;
    dff max_calc_reg_comparator_fourth_inp2_8 (.Q (\$dummy [545]), .QB (nx32319)
        , .D (nx23463), .CLK (clk)) ;
    oai21 ix23464 (.Y (nx23463), .A0 (nx32319), .A1 (nx34791), .B0 (nx32322)) ;
    oai21 ix23474 (.Y (nx23473), .A0 (nx32326), .A1 (nx34793), .B0 (nx32328)) ;
    dff max_calc_reg_comparator_fourth_inp1_8 (.Q (
        max_calc_comparator_fourth_inp1_8), .QB (nx32326), .D (nx23473), .CLK (
        clk)) ;
    oai22 ix15731 (.Y (nx15730), .A0 (nx32332), .A1 (nx32345), .B0 (
          max_calc_comparator_fourth_inp2_7), .B1 (nx32340)) ;
    oai21 ix23484 (.Y (nx23483), .A0 (nx32336), .A1 (nx34793), .B0 (nx32338)) ;
    dff max_calc_reg_comparator_fourth_inp2_7 (.Q (
        max_calc_comparator_fourth_inp2_7), .QB (nx32336), .D (nx23483), .CLK (
        clk)) ;
    nand03 ix32339 (.Y (nx32338), .A0 (label_8_output[7]), .A1 (nx35465), .A2 (
           nx34793)) ;
    dff max_calc_reg_comparator_fourth_inp1_7 (.Q (
        max_calc_comparator_fourth_inp1_7), .QB (nx32340), .D (nx23493), .CLK (
        clk)) ;
    oai21 ix23494 (.Y (nx23493), .A0 (nx32340), .A1 (nx34793), .B0 (nx32343)) ;
    nand03 ix32344 (.Y (nx32343), .A0 (label_7_output[7]), .A1 (nx35467), .A2 (
           nx34793)) ;
    aoi22 ix32346 (.Y (nx32345), .A0 (nx32347), .A1 (
          max_calc_comparator_fourth_inp1_6), .B0 (nx15536), .B1 (nx15714)) ;
    dff max_calc_reg_comparator_fourth_inp2_6 (.Q (\$dummy [546]), .QB (nx32347)
        , .D (nx23503), .CLK (clk)) ;
    oai21 ix23504 (.Y (nx23503), .A0 (nx32347), .A1 (nx34793), .B0 (nx32350)) ;
    oai21 ix23514 (.Y (nx23513), .A0 (nx32354), .A1 (nx34795), .B0 (nx32356)) ;
    dff max_calc_reg_comparator_fourth_inp1_6 (.Q (
        max_calc_comparator_fourth_inp1_6), .QB (nx32354), .D (nx23513), .CLK (
        clk)) ;
    oai22 ix15715 (.Y (nx15714), .A0 (nx32360), .A1 (nx32373), .B0 (
          max_calc_comparator_fourth_inp2_5), .B1 (nx32368)) ;
    oai21 ix23524 (.Y (nx23523), .A0 (nx32364), .A1 (nx34795), .B0 (nx32366)) ;
    dff max_calc_reg_comparator_fourth_inp2_5 (.Q (
        max_calc_comparator_fourth_inp2_5), .QB (nx32364), .D (nx23523), .CLK (
        clk)) ;
    nand03 ix32367 (.Y (nx32366), .A0 (label_8_output[5]), .A1 (nx35467), .A2 (
           nx34795)) ;
    dff max_calc_reg_comparator_fourth_inp1_5 (.Q (
        max_calc_comparator_fourth_inp1_5), .QB (nx32368), .D (nx23533), .CLK (
        clk)) ;
    oai21 ix23534 (.Y (nx23533), .A0 (nx32368), .A1 (nx34795), .B0 (nx32371)) ;
    nand03 ix32372 (.Y (nx32371), .A0 (label_7_output[5]), .A1 (nx35467), .A2 (
           nx34795)) ;
    aoi22 ix32374 (.Y (nx32373), .A0 (nx32375), .A1 (
          max_calc_comparator_fourth_inp1_4), .B0 (nx15580), .B1 (nx15698)) ;
    dff max_calc_reg_comparator_fourth_inp2_4 (.Q (\$dummy [547]), .QB (nx32375)
        , .D (nx23543), .CLK (clk)) ;
    oai21 ix23544 (.Y (nx23543), .A0 (nx32375), .A1 (nx34797), .B0 (nx32378)) ;
    oai21 ix23554 (.Y (nx23553), .A0 (nx32382), .A1 (nx34797), .B0 (nx32384)) ;
    dff max_calc_reg_comparator_fourth_inp1_4 (.Q (
        max_calc_comparator_fourth_inp1_4), .QB (nx32382), .D (nx23553), .CLK (
        clk)) ;
    oai22 ix15699 (.Y (nx15698), .A0 (nx32388), .A1 (nx32401), .B0 (
          max_calc_comparator_fourth_inp2_3), .B1 (nx32396)) ;
    oai21 ix23564 (.Y (nx23563), .A0 (nx32392), .A1 (nx34797), .B0 (nx32394)) ;
    dff max_calc_reg_comparator_fourth_inp2_3 (.Q (
        max_calc_comparator_fourth_inp2_3), .QB (nx32392), .D (nx23563), .CLK (
        clk)) ;
    nand03 ix32395 (.Y (nx32394), .A0 (label_8_output[3]), .A1 (nx35469), .A2 (
           nx34797)) ;
    dff max_calc_reg_comparator_fourth_inp1_3 (.Q (
        max_calc_comparator_fourth_inp1_3), .QB (nx32396), .D (nx23573), .CLK (
        clk)) ;
    oai21 ix23574 (.Y (nx23573), .A0 (nx32396), .A1 (nx34797), .B0 (nx32399)) ;
    nand03 ix32400 (.Y (nx32399), .A0 (label_7_output[3]), .A1 (nx35469), .A2 (
           nx34799)) ;
    aoi22 ix32402 (.Y (nx32401), .A0 (nx32403), .A1 (
          max_calc_comparator_fourth_inp1_2), .B0 (nx15624), .B1 (nx15682)) ;
    dff max_calc_reg_comparator_fourth_inp2_2 (.Q (\$dummy [548]), .QB (nx32403)
        , .D (nx23583), .CLK (clk)) ;
    oai21 ix23584 (.Y (nx23583), .A0 (nx32403), .A1 (nx34799), .B0 (nx32406)) ;
    oai21 ix23594 (.Y (nx23593), .A0 (nx32410), .A1 (nx34799), .B0 (nx32412)) ;
    dff max_calc_reg_comparator_fourth_inp1_2 (.Q (
        max_calc_comparator_fourth_inp1_2), .QB (nx32410), .D (nx23593), .CLK (
        clk)) ;
    oai21 ix15683 (.Y (nx15682), .A0 (max_calc_comparator_fourth_inp2_1), .A1 (
          nx32422), .B0 (nx32427)) ;
    oai21 ix23604 (.Y (nx23603), .A0 (nx32418), .A1 (nx34799), .B0 (nx32420)) ;
    dff max_calc_reg_comparator_fourth_inp2_1 (.Q (
        max_calc_comparator_fourth_inp2_1), .QB (nx32418), .D (nx23603), .CLK (
        clk)) ;
    nand03 ix32421 (.Y (nx32420), .A0 (label_8_output[1]), .A1 (nx35469), .A2 (
           nx34799)) ;
    dff max_calc_reg_comparator_fourth_inp1_1 (.Q (\$dummy [549]), .QB (nx32422)
        , .D (nx23613), .CLK (clk)) ;
    oai21 ix23614 (.Y (nx23613), .A0 (nx32422), .A1 (nx34801), .B0 (nx32425)) ;
    nand03 ix32426 (.Y (nx32425), .A0 (label_7_output[1]), .A1 (nx35469), .A2 (
           nx34801)) ;
    oai21 ix32428 (.Y (nx32427), .A0 (nx31429), .A1 (
          max_calc_comparator_fourth_inp1_0), .B0 (nx15646)) ;
    oai21 ix23664 (.Y (nx23663), .A0 (nx32433), .A1 (nx34801), .B0 (nx32435)) ;
    dff max_calc_reg_comparator_fourth_inp2_15 (.Q (\$dummy [550]), .QB (nx32433
        ), .D (nx23663), .CLK (clk)) ;
    nand03 ix32436 (.Y (nx32435), .A0 (label_8_output[15]), .A1 (nx35469), .A2 (
           nx34801)) ;
    dffr labelsregfile_label8_loop1_15_fx_reg_q (.Q (label_8_output[15]), .QB (
         \$dummy [551]), .D (nx23653), .CLK (clk), .R (rst)) ;
    latch lat_label_8_input_15 (.Q (label_8_input_15), .D (nx15808), .CLK (
          nx34539)) ;
    dffr reg_label_8_input_state_machine_15 (.Q (label_8_input_state_machine_15)
         , .QB (\$dummy [552]), .D (nx23643), .CLK (clk), .R (rst)) ;
    xnor2 ix15805 (.Y (nx15804), .A0 (nx15800), .A1 (nx32446)) ;
    oai22 ix15801 (.Y (nx15800), .A0 (nx31882), .A1 (nx32054), .B0 (nx32056), .B1 (
          nx31850)) ;
    oai21 ix23694 (.Y (nx23693), .A0 (nx32451), .A1 (nx34801), .B0 (nx32453)) ;
    dff max_calc_reg_comparator_fourth_inp1_15 (.Q (\$dummy [553]), .QB (nx32451
        ), .D (nx23693), .CLK (clk)) ;
    dffr labelsregfile_label7_loop1_15_fx_reg_q (.Q (label_7_output[15]), .QB (
         \$dummy [554]), .D (nx23683), .CLK (clk), .R (rst)) ;
    latch lat_label_7_input_15 (.Q (label_7_input_15), .D (nx15850), .CLK (
          nx34539)) ;
    dffr reg_label_7_input_state_machine_15 (.Q (label_7_input_state_machine_15)
         , .QB (\$dummy [555]), .D (nx23673), .CLK (clk), .R (rst)) ;
    xnor2 ix15847 (.Y (nx15846), .A0 (nx15842), .A1 (nx32464)) ;
    oai22 ix15843 (.Y (nx15842), .A0 (nx32071), .A1 (nx32243), .B0 (nx32245), .B1 (
          nx31411)) ;
    dff max_calc_reg_ans4_0 (.Q (max_calc_ans4_0), .QB (\$dummy [556]), .D (
        nx24243), .CLK (clk)) ;
    xnor2 ix17139 (.Y (nx17138), .A0 (nx32470), .A1 (nx17136)) ;
    aoi22 ix32471 (.Y (nx32470), .A0 (nx32472), .A1 (
          max_calc_comparator_second_inp1_14), .B0 (nx15908), .B1 (nx17054)) ;
    dff max_calc_reg_comparator_second_inp2_14 (.Q (\$dummy [557]), .QB (nx32472
        ), .D (nx23713), .CLK (clk)) ;
    oai21 ix23714 (.Y (nx23713), .A0 (nx32472), .A1 (nx34803), .B0 (nx32475)) ;
    nand03 ix32476 (.Y (nx32475), .A0 (nx35175), .A1 (nx15896), .A2 (nx34803)) ;
    dffr labelsregfile_label4_loop1_14_fx_reg_q (.Q (label_4_output[14]), .QB (
         nx32660), .D (nx14953), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_14 (.Q (label_4_input_14), .D (nx2186), .CLK (
          nx34543)) ;
    dffr reg_label_4_input_state_machine_14 (.Q (label_4_input_state_machine_14)
         , .QB (\$dummy [558]), .D (nx14943), .CLK (clk), .R (rst)) ;
    xor2 ix2183 (.Y (nx2182), .A0 (nx32486), .A1 (nx32658)) ;
    aoi22 ix32487 (.Y (nx32486), .A0 (label_4_output[13]), .A1 (
          booth_booth_integration_output_3_13), .B0 (nx2140), .B1 (nx12959)) ;
    dffr labelsregfile_label4_loop1_13_fx_reg_q (.Q (label_4_output[13]), .QB (
         \$dummy [559]), .D (nx14933), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_13 (.Q (label_4_input_13), .D (nx2154), .CLK (
          nx34543)) ;
    dffr reg_label_4_input_state_machine_13 (.Q (label_4_input_state_machine_13)
         , .QB (\$dummy [560]), .D (nx14923), .CLK (clk), .R (rst)) ;
    xnor2 ix2151 (.Y (nx2150), .A0 (nx2140), .A1 (nx32654)) ;
    oai22 ix2141 (.Y (nx2140), .A0 (nx32497), .A1 (nx32643), .B0 (nx32653), .B1 (
          nx30970)) ;
    aoi22 ix32498 (.Y (nx32497), .A0 (label_4_output[11]), .A1 (
          booth_booth_integration_output_3_11), .B0 (nx2076), .B1 (nx12955)) ;
    dffr labelsregfile_label4_loop1_11_fx_reg_q (.Q (label_4_output[11]), .QB (
         \$dummy [561]), .D (nx14893), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_11 (.Q (label_4_input_11), .D (nx2090), .CLK (
          nx34541)) ;
    dffr reg_label_4_input_state_machine_11 (.Q (label_4_input_state_machine_11)
         , .QB (\$dummy [562]), .D (nx14883), .CLK (clk), .R (rst)) ;
    xnor2 ix2087 (.Y (nx2086), .A0 (nx2076), .A1 (nx32639)) ;
    oai22 ix2077 (.Y (nx2076), .A0 (nx32508), .A1 (nx32628), .B0 (nx32638), .B1 (
          nx30972)) ;
    aoi22 ix32509 (.Y (nx32508), .A0 (label_4_output[9]), .A1 (
          booth_booth_integration_output_3_9), .B0 (nx2012), .B1 (nx12953)) ;
    dffr labelsregfile_label4_loop1_9_fx_reg_q (.Q (label_4_output[9]), .QB (
         \$dummy [563]), .D (nx14853), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_9 (.Q (label_4_input_9), .D (nx2026), .CLK (nx34541)
          ) ;
    dffr reg_label_4_input_state_machine_9 (.Q (label_4_input_state_machine_9), 
         .QB (\$dummy [564]), .D (nx14843), .CLK (clk), .R (rst)) ;
    xnor2 ix2023 (.Y (nx2022), .A0 (nx2012), .A1 (nx32624)) ;
    oai22 ix2013 (.Y (nx2012), .A0 (nx32519), .A1 (nx32613), .B0 (nx32623), .B1 (
          nx30974)) ;
    aoi22 ix32520 (.Y (nx32519), .A0 (label_4_output[7]), .A1 (
          booth_booth_integration_output_3_7), .B0 (nx1948), .B1 (nx12949)) ;
    dffr labelsregfile_label4_loop1_7_fx_reg_q (.Q (label_4_output[7]), .QB (
         \$dummy [565]), .D (nx14813), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_7 (.Q (label_4_input_7), .D (nx1962), .CLK (nx34541)
          ) ;
    dffr reg_label_4_input_state_machine_7 (.Q (label_4_input_state_machine_7), 
         .QB (\$dummy [566]), .D (nx14803), .CLK (clk), .R (rst)) ;
    xnor2 ix1959 (.Y (nx1958), .A0 (nx1948), .A1 (nx32609)) ;
    oai22 ix1949 (.Y (nx1948), .A0 (nx32530), .A1 (nx32598), .B0 (nx32608), .B1 (
          nx30976)) ;
    aoi22 ix32531 (.Y (nx32530), .A0 (label_4_output[5]), .A1 (
          booth_booth_integration_output_3_5), .B0 (nx1884), .B1 (nx12946)) ;
    dffr labelsregfile_label4_loop1_5_fx_reg_q (.Q (label_4_output[5]), .QB (
         \$dummy [567]), .D (nx14773), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_5 (.Q (label_4_input_5), .D (nx1898), .CLK (nx34539)
          ) ;
    dffr reg_label_4_input_state_machine_5 (.Q (label_4_input_state_machine_5), 
         .QB (\$dummy [568]), .D (nx14763), .CLK (clk), .R (rst)) ;
    xnor2 ix1895 (.Y (nx1894), .A0 (nx1884), .A1 (nx32594)) ;
    oai22 ix1885 (.Y (nx1884), .A0 (nx32541), .A1 (nx32583), .B0 (nx32593), .B1 (
          nx30978)) ;
    aoi22 ix32542 (.Y (nx32541), .A0 (label_4_output[3]), .A1 (
          booth_booth_integration_output_3_3), .B0 (nx1820), .B1 (nx12943)) ;
    dffr labelsregfile_label4_loop1_3_fx_reg_q (.Q (label_4_output[3]), .QB (
         \$dummy [569]), .D (nx14733), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_3 (.Q (label_4_input_3), .D (nx1834), .CLK (nx34539)
          ) ;
    dffr reg_label_4_input_state_machine_3 (.Q (label_4_input_state_machine_3), 
         .QB (\$dummy [570]), .D (nx14723), .CLK (clk), .R (rst)) ;
    xnor2 ix1831 (.Y (nx1830), .A0 (nx1820), .A1 (nx32579)) ;
    oai22 ix1821 (.Y (nx1820), .A0 (nx32552), .A1 (nx32568), .B0 (nx32578), .B1 (
          nx30980)) ;
    aoi32 ix32553 (.Y (nx32552), .A0 (label_4_output[0]), .A1 (nx35719), .A2 (
          nx12939), .B0 (label_4_output[1]), .B1 (
          booth_booth_integration_output_3_1)) ;
    dffr labelsregfile_label4_loop1_1_fx_reg_q (.Q (label_4_output[1]), .QB (
         \$dummy [571]), .D (nx14693), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_1 (.Q (label_4_input_1), .D (nx1770), .CLK (nx34539)
          ) ;
    dffr reg_label_4_input_state_machine_1 (.Q (label_4_input_state_machine_1), 
         .QB (\$dummy [572]), .D (nx14683), .CLK (clk), .R (rst)) ;
    xor2 ix1767 (.Y (nx1766), .A0 (nx32563), .A1 (nx32565)) ;
    nand02 ix32564 (.Y (nx32563), .A0 (label_4_output[0]), .A1 (nx35719)) ;
    xnor2 ix32566 (.Y (nx32565), .A0 (booth_booth_integration_output_3_1), .A1 (
          label_4_output[1])) ;
    dffr labelsregfile_label4_loop1_2_fx_reg_q (.Q (label_4_output[2]), .QB (
         nx32578), .D (nx14713), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_2 (.Q (label_4_input_2), .D (nx1802), .CLK (nx34539)
          ) ;
    dffr reg_label_4_input_state_machine_2 (.Q (label_4_input_state_machine_2), 
         .QB (\$dummy [573]), .D (nx14703), .CLK (clk), .R (rst)) ;
    xor2 ix1799 (.Y (nx1798), .A0 (nx32552), .A1 (nx32568)) ;
    xnor2 ix32580 (.Y (nx32579), .A0 (booth_booth_integration_output_3_3), .A1 (
          label_4_output[3])) ;
    dffr labelsregfile_label4_loop1_4_fx_reg_q (.Q (label_4_output[4]), .QB (
         nx32593), .D (nx14753), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_4 (.Q (label_4_input_4), .D (nx1866), .CLK (nx34539)
          ) ;
    dffr reg_label_4_input_state_machine_4 (.Q (label_4_input_state_machine_4), 
         .QB (\$dummy [574]), .D (nx14743), .CLK (clk), .R (rst)) ;
    xor2 ix1863 (.Y (nx1862), .A0 (nx32541), .A1 (nx32583)) ;
    xnor2 ix32595 (.Y (nx32594), .A0 (booth_booth_integration_output_3_5), .A1 (
          label_4_output[5])) ;
    dffr labelsregfile_label4_loop1_6_fx_reg_q (.Q (label_4_output[6]), .QB (
         nx32608), .D (nx14793), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_6 (.Q (label_4_input_6), .D (nx1930), .CLK (nx34541)
          ) ;
    dffr reg_label_4_input_state_machine_6 (.Q (label_4_input_state_machine_6), 
         .QB (\$dummy [575]), .D (nx14783), .CLK (clk), .R (rst)) ;
    xor2 ix1927 (.Y (nx1926), .A0 (nx32530), .A1 (nx32598)) ;
    xnor2 ix32610 (.Y (nx32609), .A0 (booth_booth_integration_output_3_7), .A1 (
          label_4_output[7])) ;
    dffr labelsregfile_label4_loop1_8_fx_reg_q (.Q (label_4_output[8]), .QB (
         nx32623), .D (nx14833), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_8 (.Q (label_4_input_8), .D (nx1994), .CLK (nx34541)
          ) ;
    dffr reg_label_4_input_state_machine_8 (.Q (label_4_input_state_machine_8), 
         .QB (\$dummy [576]), .D (nx14823), .CLK (clk), .R (rst)) ;
    xor2 ix1991 (.Y (nx1990), .A0 (nx32519), .A1 (nx32613)) ;
    xnor2 ix32625 (.Y (nx32624), .A0 (booth_booth_integration_output_3_9), .A1 (
          label_4_output[9])) ;
    dffr labelsregfile_label4_loop1_10_fx_reg_q (.Q (label_4_output[10]), .QB (
         nx32638), .D (nx14873), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_10 (.Q (label_4_input_10), .D (nx2058), .CLK (
          nx34541)) ;
    dffr reg_label_4_input_state_machine_10 (.Q (label_4_input_state_machine_10)
         , .QB (\$dummy [577]), .D (nx14863), .CLK (clk), .R (rst)) ;
    xor2 ix2055 (.Y (nx2054), .A0 (nx32508), .A1 (nx32628)) ;
    xnor2 ix32640 (.Y (nx32639), .A0 (booth_booth_integration_output_3_11), .A1 (
          label_4_output[11])) ;
    dffr labelsregfile_label4_loop1_12_fx_reg_q (.Q (label_4_output[12]), .QB (
         nx32653), .D (nx14913), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_12 (.Q (label_4_input_12), .D (nx2122), .CLK (
          nx34541)) ;
    dffr reg_label_4_input_state_machine_12 (.Q (label_4_input_state_machine_12)
         , .QB (\$dummy [578]), .D (nx14903), .CLK (clk), .R (rst)) ;
    xor2 ix2119 (.Y (nx2118), .A0 (nx32497), .A1 (nx32643)) ;
    xnor2 ix32655 (.Y (nx32654), .A0 (booth_booth_integration_output_3_13), .A1 (
          label_4_output[13])) ;
    dff max_calc_reg_ans4_14 (.Q (max_calc_ans4_14), .QB (nx32665), .D (nx23703)
        , .CLK (clk)) ;
    oai21 ix21674 (.Y (nx21673), .A0 (nx32669), .A1 (nx34803), .B0 (nx32671)) ;
    dff max_calc_reg_comparator_second_inp1_14 (.Q (
        max_calc_comparator_second_inp1_14), .QB (nx32669), .D (nx21673), .CLK (
        clk)) ;
    nand03 ix32672 (.Y (nx32671), .A0 (nx35175), .A1 (nx12712), .A2 (nx34803)) ;
    dffr labelsregfile_label3_loop1_14_fx_reg_q (.Q (label_3_output[14]), .QB (
         nx32856), .D (nx15803), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_14 (.Q (label_3_input_14), .D (nx3524), .CLK (
          nx34547)) ;
    dffr reg_label_3_input_state_machine_14 (.Q (label_3_input_state_machine_14)
         , .QB (\$dummy [579]), .D (nx15793), .CLK (clk), .R (rst)) ;
    xor2 ix3521 (.Y (nx3520), .A0 (nx32682), .A1 (nx32854)) ;
    aoi22 ix32683 (.Y (nx32682), .A0 (label_3_output[13]), .A1 (
          booth_booth_integration_output_2_13), .B0 (nx3478), .B1 (nx13011)) ;
    dffr labelsregfile_label3_loop1_13_fx_reg_q (.Q (label_3_output[13]), .QB (
         \$dummy [580]), .D (nx15783), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_13 (.Q (label_3_input_13), .D (nx3492), .CLK (
          nx34547)) ;
    dffr reg_label_3_input_state_machine_13 (.Q (label_3_input_state_machine_13)
         , .QB (\$dummy [581]), .D (nx15773), .CLK (clk), .R (rst)) ;
    xnor2 ix3489 (.Y (nx3488), .A0 (nx3478), .A1 (nx32850)) ;
    oai22 ix3479 (.Y (nx3478), .A0 (nx32693), .A1 (nx32839), .B0 (nx32849), .B1 (
          nx29041)) ;
    aoi22 ix32694 (.Y (nx32693), .A0 (label_3_output[11]), .A1 (
          booth_booth_integration_output_2_11), .B0 (nx3414), .B1 (nx13007)) ;
    dffr labelsregfile_label3_loop1_11_fx_reg_q (.Q (label_3_output[11]), .QB (
         \$dummy [582]), .D (nx15743), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_11 (.Q (label_3_input_11), .D (nx3428), .CLK (
          nx34545)) ;
    dffr reg_label_3_input_state_machine_11 (.Q (label_3_input_state_machine_11)
         , .QB (\$dummy [583]), .D (nx15733), .CLK (clk), .R (rst)) ;
    xnor2 ix3425 (.Y (nx3424), .A0 (nx3414), .A1 (nx32835)) ;
    oai22 ix3415 (.Y (nx3414), .A0 (nx32704), .A1 (nx32824), .B0 (nx32834), .B1 (
          nx29043)) ;
    aoi22 ix32705 (.Y (nx32704), .A0 (label_3_output[9]), .A1 (
          booth_booth_integration_output_2_9), .B0 (nx3350), .B1 (nx13003)) ;
    dffr labelsregfile_label3_loop1_9_fx_reg_q (.Q (label_3_output[9]), .QB (
         \$dummy [584]), .D (nx15703), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_9 (.Q (label_3_input_9), .D (nx3364), .CLK (nx34545)
          ) ;
    dffr reg_label_3_input_state_machine_9 (.Q (label_3_input_state_machine_9), 
         .QB (\$dummy [585]), .D (nx15693), .CLK (clk), .R (rst)) ;
    xnor2 ix3361 (.Y (nx3360), .A0 (nx3350), .A1 (nx32820)) ;
    oai22 ix3351 (.Y (nx3350), .A0 (nx32715), .A1 (nx32809), .B0 (nx32819), .B1 (
          nx29045)) ;
    aoi22 ix32716 (.Y (nx32715), .A0 (label_3_output[7]), .A1 (
          booth_booth_integration_output_2_7), .B0 (nx3286), .B1 (nx13001)) ;
    dffr labelsregfile_label3_loop1_7_fx_reg_q (.Q (label_3_output[7]), .QB (
         \$dummy [586]), .D (nx15663), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_7 (.Q (label_3_input_7), .D (nx3300), .CLK (nx34545)
          ) ;
    dffr reg_label_3_input_state_machine_7 (.Q (label_3_input_state_machine_7), 
         .QB (\$dummy [587]), .D (nx15653), .CLK (clk), .R (rst)) ;
    xnor2 ix3297 (.Y (nx3296), .A0 (nx3286), .A1 (nx32805)) ;
    oai22 ix3287 (.Y (nx3286), .A0 (nx32726), .A1 (nx32794), .B0 (nx32804), .B1 (
          nx29047)) ;
    aoi22 ix32727 (.Y (nx32726), .A0 (label_3_output[5]), .A1 (
          booth_booth_integration_output_2_5), .B0 (nx3222), .B1 (nx12997)) ;
    dffr labelsregfile_label3_loop1_5_fx_reg_q (.Q (label_3_output[5]), .QB (
         \$dummy [588]), .D (nx15623), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_5 (.Q (label_3_input_5), .D (nx3236), .CLK (nx34543)
          ) ;
    dffr reg_label_3_input_state_machine_5 (.Q (label_3_input_state_machine_5), 
         .QB (\$dummy [589]), .D (nx15613), .CLK (clk), .R (rst)) ;
    xnor2 ix3233 (.Y (nx3232), .A0 (nx3222), .A1 (nx32790)) ;
    oai22 ix3223 (.Y (nx3222), .A0 (nx32737), .A1 (nx32779), .B0 (nx32789), .B1 (
          nx29049)) ;
    aoi22 ix32738 (.Y (nx32737), .A0 (label_3_output[3]), .A1 (
          booth_booth_integration_output_2_3), .B0 (nx3158), .B1 (nx12994)) ;
    dffr labelsregfile_label3_loop1_3_fx_reg_q (.Q (label_3_output[3]), .QB (
         \$dummy [590]), .D (nx15583), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_3 (.Q (label_3_input_3), .D (nx3172), .CLK (nx34543)
          ) ;
    dffr reg_label_3_input_state_machine_3 (.Q (label_3_input_state_machine_3), 
         .QB (\$dummy [591]), .D (nx15573), .CLK (clk), .R (rst)) ;
    xnor2 ix3169 (.Y (nx3168), .A0 (nx3158), .A1 (nx32775)) ;
    oai22 ix3159 (.Y (nx3158), .A0 (nx32748), .A1 (nx32764), .B0 (nx32774), .B1 (
          nx29051)) ;
    aoi32 ix32749 (.Y (nx32748), .A0 (label_3_output[0]), .A1 (nx35723), .A2 (
          nx12991), .B0 (label_3_output[1]), .B1 (
          booth_booth_integration_output_2_1)) ;
    dffr labelsregfile_label3_loop1_1_fx_reg_q (.Q (label_3_output[1]), .QB (
         \$dummy [592]), .D (nx15543), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_1 (.Q (label_3_input_1), .D (nx3108), .CLK (nx34543)
          ) ;
    dffr reg_label_3_input_state_machine_1 (.Q (label_3_input_state_machine_1), 
         .QB (\$dummy [593]), .D (nx15533), .CLK (clk), .R (rst)) ;
    xor2 ix3105 (.Y (nx3104), .A0 (nx32759), .A1 (nx32761)) ;
    nand02 ix32760 (.Y (nx32759), .A0 (label_3_output[0]), .A1 (nx35723)) ;
    xnor2 ix32762 (.Y (nx32761), .A0 (booth_booth_integration_output_2_1), .A1 (
          label_3_output[1])) ;
    dffr labelsregfile_label3_loop1_2_fx_reg_q (.Q (label_3_output[2]), .QB (
         nx32774), .D (nx15563), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_2 (.Q (label_3_input_2), .D (nx3140), .CLK (nx34543)
          ) ;
    dffr reg_label_3_input_state_machine_2 (.Q (label_3_input_state_machine_2), 
         .QB (\$dummy [594]), .D (nx15553), .CLK (clk), .R (rst)) ;
    xor2 ix3137 (.Y (nx3136), .A0 (nx32748), .A1 (nx32764)) ;
    xnor2 ix32776 (.Y (nx32775), .A0 (booth_booth_integration_output_2_3), .A1 (
          label_3_output[3])) ;
    dffr labelsregfile_label3_loop1_4_fx_reg_q (.Q (label_3_output[4]), .QB (
         nx32789), .D (nx15603), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_4 (.Q (label_3_input_4), .D (nx3204), .CLK (nx34543)
          ) ;
    dffr reg_label_3_input_state_machine_4 (.Q (label_3_input_state_machine_4), 
         .QB (\$dummy [595]), .D (nx15593), .CLK (clk), .R (rst)) ;
    xor2 ix3201 (.Y (nx3200), .A0 (nx32737), .A1 (nx32779)) ;
    xnor2 ix32791 (.Y (nx32790), .A0 (booth_booth_integration_output_2_5), .A1 (
          label_3_output[5])) ;
    dffr labelsregfile_label3_loop1_6_fx_reg_q (.Q (label_3_output[6]), .QB (
         nx32804), .D (nx15643), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_6 (.Q (label_3_input_6), .D (nx3268), .CLK (nx34545)
          ) ;
    dffr reg_label_3_input_state_machine_6 (.Q (label_3_input_state_machine_6), 
         .QB (\$dummy [596]), .D (nx15633), .CLK (clk), .R (rst)) ;
    xor2 ix3265 (.Y (nx3264), .A0 (nx32726), .A1 (nx32794)) ;
    xnor2 ix32806 (.Y (nx32805), .A0 (booth_booth_integration_output_2_7), .A1 (
          label_3_output[7])) ;
    dffr labelsregfile_label3_loop1_8_fx_reg_q (.Q (label_3_output[8]), .QB (
         nx32819), .D (nx15683), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_8 (.Q (label_3_input_8), .D (nx3332), .CLK (nx34545)
          ) ;
    dffr reg_label_3_input_state_machine_8 (.Q (label_3_input_state_machine_8), 
         .QB (\$dummy [597]), .D (nx15673), .CLK (clk), .R (rst)) ;
    xor2 ix3329 (.Y (nx3328), .A0 (nx32715), .A1 (nx32809)) ;
    xnor2 ix32821 (.Y (nx32820), .A0 (booth_booth_integration_output_2_9), .A1 (
          label_3_output[9])) ;
    dffr labelsregfile_label3_loop1_10_fx_reg_q (.Q (label_3_output[10]), .QB (
         nx32834), .D (nx15723), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_10 (.Q (label_3_input_10), .D (nx3396), .CLK (
          nx34545)) ;
    dffr reg_label_3_input_state_machine_10 (.Q (label_3_input_state_machine_10)
         , .QB (\$dummy [598]), .D (nx15713), .CLK (clk), .R (rst)) ;
    xor2 ix3393 (.Y (nx3392), .A0 (nx32704), .A1 (nx32824)) ;
    xnor2 ix32836 (.Y (nx32835), .A0 (booth_booth_integration_output_2_11), .A1 (
          label_3_output[11])) ;
    dffr labelsregfile_label3_loop1_12_fx_reg_q (.Q (label_3_output[12]), .QB (
         nx32849), .D (nx15763), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_12 (.Q (label_3_input_12), .D (nx3460), .CLK (
          nx34545)) ;
    dffr reg_label_3_input_state_machine_12 (.Q (label_3_input_state_machine_12)
         , .QB (\$dummy [599]), .D (nx15753), .CLK (clk), .R (rst)) ;
    xor2 ix3457 (.Y (nx3456), .A0 (nx32693), .A1 (nx32839)) ;
    xnor2 ix32851 (.Y (nx32850), .A0 (booth_booth_integration_output_2_13), .A1 (
          label_3_output[13])) ;
    dff max_calc_reg_ans3_14 (.Q (max_calc_ans3_14), .QB (nx32861), .D (nx21663)
        , .CLK (clk)) ;
    oai22 ix17055 (.Y (nx17054), .A0 (nx32865), .A1 (nx32892), .B0 (
          max_calc_comparator_second_inp2_13), .B1 (nx32880)) ;
    oai21 ix23734 (.Y (nx23733), .A0 (nx32869), .A1 (nx34803), .B0 (nx32871)) ;
    dff max_calc_reg_comparator_second_inp2_13 (.Q (
        max_calc_comparator_second_inp2_13), .QB (nx32869), .D (nx23733), .CLK (
        clk)) ;
    nand03 ix32872 (.Y (nx32871), .A0 (nx35175), .A1 (nx15934), .A2 (nx34803)) ;
    dff max_calc_reg_ans4_13 (.Q (max_calc_ans4_13), .QB (\$dummy [600]), .D (
        nx23723), .CLK (clk)) ;
    dff max_calc_reg_comparator_second_inp1_13 (.Q (
        max_calc_comparator_second_inp1_13), .QB (nx32880), .D (nx23753), .CLK (
        clk)) ;
    oai21 ix23754 (.Y (nx23753), .A0 (nx32880), .A1 (nx34803), .B0 (nx32883)) ;
    nand03 ix32884 (.Y (nx32883), .A0 (nx35175), .A1 (nx15970), .A2 (nx34805)) ;
    dff max_calc_reg_ans3_13 (.Q (max_calc_ans3_13), .QB (\$dummy [601]), .D (
        nx23743), .CLK (clk)) ;
    aoi22 ix32893 (.Y (nx32892), .A0 (nx32894), .A1 (
          max_calc_comparator_second_inp1_12), .B0 (nx16056), .B1 (nx17038)) ;
    dff max_calc_reg_comparator_second_inp2_12 (.Q (\$dummy [602]), .QB (nx32894
        ), .D (nx23773), .CLK (clk)) ;
    oai21 ix23774 (.Y (nx23773), .A0 (nx32894), .A1 (nx34805), .B0 (nx32897)) ;
    nand03 ix32898 (.Y (nx32897), .A0 (nx35175), .A1 (nx16008), .A2 (nx34805)) ;
    dff max_calc_reg_ans4_12 (.Q (max_calc_ans4_12), .QB (nx32904), .D (nx23763)
        , .CLK (clk)) ;
    oai21 ix23794 (.Y (nx23793), .A0 (nx32908), .A1 (nx34805), .B0 (nx32910)) ;
    dff max_calc_reg_comparator_second_inp1_12 (.Q (
        max_calc_comparator_second_inp1_12), .QB (nx32908), .D (nx23793), .CLK (
        clk)) ;
    nand03 ix32911 (.Y (nx32910), .A0 (nx35175), .A1 (nx16044), .A2 (nx34805)) ;
    dff max_calc_reg_ans3_12 (.Q (max_calc_ans3_12), .QB (nx32917), .D (nx23783)
        , .CLK (clk)) ;
    oai22 ix17039 (.Y (nx17038), .A0 (nx32921), .A1 (nx32948), .B0 (
          max_calc_comparator_second_inp2_11), .B1 (nx32936)) ;
    oai21 ix23814 (.Y (nx23813), .A0 (nx32925), .A1 (nx34805), .B0 (nx32927)) ;
    dff max_calc_reg_comparator_second_inp2_11 (.Q (
        max_calc_comparator_second_inp2_11), .QB (nx32925), .D (nx23813), .CLK (
        clk)) ;
    nand03 ix32928 (.Y (nx32927), .A0 (nx35177), .A1 (nx16082), .A2 (nx34805)) ;
    dff max_calc_reg_ans4_11 (.Q (max_calc_ans4_11), .QB (\$dummy [603]), .D (
        nx23803), .CLK (clk)) ;
    dff max_calc_reg_comparator_second_inp1_11 (.Q (
        max_calc_comparator_second_inp1_11), .QB (nx32936), .D (nx23833), .CLK (
        clk)) ;
    oai21 ix23834 (.Y (nx23833), .A0 (nx32936), .A1 (nx34807), .B0 (nx32939)) ;
    nand03 ix32940 (.Y (nx32939), .A0 (nx35177), .A1 (nx16118), .A2 (nx34807)) ;
    dff max_calc_reg_ans3_11 (.Q (max_calc_ans3_11), .QB (\$dummy [604]), .D (
        nx23823), .CLK (clk)) ;
    aoi22 ix32949 (.Y (nx32948), .A0 (nx32950), .A1 (
          max_calc_comparator_second_inp1_10), .B0 (nx16204), .B1 (nx17022)) ;
    dff max_calc_reg_comparator_second_inp2_10 (.Q (\$dummy [605]), .QB (nx32950
        ), .D (nx23853), .CLK (clk)) ;
    oai21 ix23854 (.Y (nx23853), .A0 (nx32950), .A1 (nx34807), .B0 (nx32953)) ;
    nand03 ix32954 (.Y (nx32953), .A0 (nx35177), .A1 (nx16156), .A2 (nx34807)) ;
    dff max_calc_reg_ans4_10 (.Q (max_calc_ans4_10), .QB (nx32960), .D (nx23843)
        , .CLK (clk)) ;
    oai21 ix23874 (.Y (nx23873), .A0 (nx32964), .A1 (nx34807), .B0 (nx32966)) ;
    dff max_calc_reg_comparator_second_inp1_10 (.Q (
        max_calc_comparator_second_inp1_10), .QB (nx32964), .D (nx23873), .CLK (
        clk)) ;
    nand03 ix32967 (.Y (nx32966), .A0 (nx35177), .A1 (nx16192), .A2 (nx34807)) ;
    dff max_calc_reg_ans3_10 (.Q (max_calc_ans3_10), .QB (nx32973), .D (nx23863)
        , .CLK (clk)) ;
    oai22 ix17023 (.Y (nx17022), .A0 (nx32977), .A1 (nx33004), .B0 (
          max_calc_comparator_second_inp2_9), .B1 (nx32992)) ;
    oai21 ix23894 (.Y (nx23893), .A0 (nx32981), .A1 (nx34807), .B0 (nx32983)) ;
    dff max_calc_reg_comparator_second_inp2_9 (.Q (
        max_calc_comparator_second_inp2_9), .QB (nx32981), .D (nx23893), .CLK (
        clk)) ;
    nand03 ix32984 (.Y (nx32983), .A0 (nx35177), .A1 (nx16230), .A2 (nx34809)) ;
    dff max_calc_reg_ans4_9 (.Q (max_calc_ans4_9), .QB (\$dummy [606]), .D (
        nx23883), .CLK (clk)) ;
    dff max_calc_reg_comparator_second_inp1_9 (.Q (
        max_calc_comparator_second_inp1_9), .QB (nx32992), .D (nx23913), .CLK (
        clk)) ;
    oai21 ix23914 (.Y (nx23913), .A0 (nx32992), .A1 (nx34809), .B0 (nx32995)) ;
    nand03 ix32996 (.Y (nx32995), .A0 (nx35177), .A1 (nx16266), .A2 (nx34809)) ;
    dff max_calc_reg_ans3_9 (.Q (max_calc_ans3_9), .QB (\$dummy [607]), .D (
        nx23903), .CLK (clk)) ;
    aoi22 ix33005 (.Y (nx33004), .A0 (nx33006), .A1 (
          max_calc_comparator_second_inp1_8), .B0 (nx16352), .B1 (nx17006)) ;
    dff max_calc_reg_comparator_second_inp2_8 (.Q (\$dummy [608]), .QB (nx33006)
        , .D (nx23933), .CLK (clk)) ;
    oai21 ix23934 (.Y (nx23933), .A0 (nx33006), .A1 (nx34809), .B0 (nx33009)) ;
    nand03 ix33010 (.Y (nx33009), .A0 (nx35177), .A1 (nx16304), .A2 (nx34809)) ;
    dff max_calc_reg_ans4_8 (.Q (max_calc_ans4_8), .QB (nx33016), .D (nx23923), 
        .CLK (clk)) ;
    oai21 ix23954 (.Y (nx23953), .A0 (nx33020), .A1 (nx34809), .B0 (nx33022)) ;
    dff max_calc_reg_comparator_second_inp1_8 (.Q (
        max_calc_comparator_second_inp1_8), .QB (nx33020), .D (nx23953), .CLK (
        clk)) ;
    nand03 ix33023 (.Y (nx33022), .A0 (nx35179), .A1 (nx16340), .A2 (nx34809)) ;
    dff max_calc_reg_ans3_8 (.Q (max_calc_ans3_8), .QB (nx33029), .D (nx23943), 
        .CLK (clk)) ;
    oai22 ix17007 (.Y (nx17006), .A0 (nx33033), .A1 (nx33060), .B0 (
          max_calc_comparator_second_inp2_7), .B1 (nx33048)) ;
    oai21 ix23974 (.Y (nx23973), .A0 (nx33037), .A1 (nx34811), .B0 (nx33039)) ;
    dff max_calc_reg_comparator_second_inp2_7 (.Q (
        max_calc_comparator_second_inp2_7), .QB (nx33037), .D (nx23973), .CLK (
        clk)) ;
    nand03 ix33040 (.Y (nx33039), .A0 (nx35179), .A1 (nx16378), .A2 (nx34811)) ;
    dff max_calc_reg_ans4_7 (.Q (max_calc_ans4_7), .QB (\$dummy [609]), .D (
        nx23963), .CLK (clk)) ;
    dff max_calc_reg_comparator_second_inp1_7 (.Q (
        max_calc_comparator_second_inp1_7), .QB (nx33048), .D (nx23993), .CLK (
        clk)) ;
    oai21 ix23994 (.Y (nx23993), .A0 (nx33048), .A1 (nx34811), .B0 (nx33051)) ;
    nand03 ix33052 (.Y (nx33051), .A0 (nx35179), .A1 (nx16414), .A2 (nx34811)) ;
    dff max_calc_reg_ans3_7 (.Q (max_calc_ans3_7), .QB (\$dummy [610]), .D (
        nx23983), .CLK (clk)) ;
    aoi22 ix33061 (.Y (nx33060), .A0 (nx33062), .A1 (
          max_calc_comparator_second_inp1_6), .B0 (nx16500), .B1 (nx16990)) ;
    dff max_calc_reg_comparator_second_inp2_6 (.Q (\$dummy [611]), .QB (nx33062)
        , .D (nx24013), .CLK (clk)) ;
    oai21 ix24014 (.Y (nx24013), .A0 (nx33062), .A1 (nx34811), .B0 (nx33065)) ;
    nand03 ix33066 (.Y (nx33065), .A0 (nx35179), .A1 (nx16452), .A2 (nx34811)) ;
    dff max_calc_reg_ans4_6 (.Q (max_calc_ans4_6), .QB (nx33072), .D (nx24003), 
        .CLK (clk)) ;
    oai21 ix24034 (.Y (nx24033), .A0 (nx33076), .A1 (nx34811), .B0 (nx33078)) ;
    dff max_calc_reg_comparator_second_inp1_6 (.Q (
        max_calc_comparator_second_inp1_6), .QB (nx33076), .D (nx24033), .CLK (
        clk)) ;
    nand03 ix33079 (.Y (nx33078), .A0 (nx35179), .A1 (nx16488), .A2 (nx34813)) ;
    dff max_calc_reg_ans3_6 (.Q (max_calc_ans3_6), .QB (nx33085), .D (nx24023), 
        .CLK (clk)) ;
    oai22 ix16991 (.Y (nx16990), .A0 (nx33089), .A1 (nx33116), .B0 (
          max_calc_comparator_second_inp2_5), .B1 (nx33104)) ;
    oai21 ix24054 (.Y (nx24053), .A0 (nx33093), .A1 (nx34813), .B0 (nx33095)) ;
    dff max_calc_reg_comparator_second_inp2_5 (.Q (
        max_calc_comparator_second_inp2_5), .QB (nx33093), .D (nx24053), .CLK (
        clk)) ;
    nand03 ix33096 (.Y (nx33095), .A0 (nx35179), .A1 (nx16526), .A2 (nx34813)) ;
    dff max_calc_reg_ans4_5 (.Q (max_calc_ans4_5), .QB (\$dummy [612]), .D (
        nx24043), .CLK (clk)) ;
    dff max_calc_reg_comparator_second_inp1_5 (.Q (
        max_calc_comparator_second_inp1_5), .QB (nx33104), .D (nx24073), .CLK (
        clk)) ;
    oai21 ix24074 (.Y (nx24073), .A0 (nx33104), .A1 (nx34813), .B0 (nx33107)) ;
    nand03 ix33108 (.Y (nx33107), .A0 (nx35179), .A1 (nx16562), .A2 (nx34813)) ;
    dff max_calc_reg_ans3_5 (.Q (max_calc_ans3_5), .QB (\$dummy [613]), .D (
        nx24063), .CLK (clk)) ;
    aoi22 ix33117 (.Y (nx33116), .A0 (nx33118), .A1 (
          max_calc_comparator_second_inp1_4), .B0 (nx16648), .B1 (nx16974)) ;
    dff max_calc_reg_comparator_second_inp2_4 (.Q (\$dummy [614]), .QB (nx33118)
        , .D (nx24093), .CLK (clk)) ;
    oai21 ix24094 (.Y (nx24093), .A0 (nx33118), .A1 (nx34813), .B0 (nx33121)) ;
    nand03 ix33122 (.Y (nx33121), .A0 (nx35181), .A1 (nx16600), .A2 (nx34813)) ;
    dff max_calc_reg_ans4_4 (.Q (max_calc_ans4_4), .QB (nx33128), .D (nx24083), 
        .CLK (clk)) ;
    oai21 ix24114 (.Y (nx24113), .A0 (nx33132), .A1 (nx34815), .B0 (nx33134)) ;
    dff max_calc_reg_comparator_second_inp1_4 (.Q (
        max_calc_comparator_second_inp1_4), .QB (nx33132), .D (nx24113), .CLK (
        clk)) ;
    nand03 ix33135 (.Y (nx33134), .A0 (nx35181), .A1 (nx16636), .A2 (nx34815)) ;
    dff max_calc_reg_ans3_4 (.Q (max_calc_ans3_4), .QB (nx33141), .D (nx24103), 
        .CLK (clk)) ;
    oai22 ix16975 (.Y (nx16974), .A0 (nx33145), .A1 (nx33172), .B0 (
          max_calc_comparator_second_inp2_3), .B1 (nx33160)) ;
    oai21 ix24134 (.Y (nx24133), .A0 (nx33149), .A1 (nx34815), .B0 (nx33151)) ;
    dff max_calc_reg_comparator_second_inp2_3 (.Q (
        max_calc_comparator_second_inp2_3), .QB (nx33149), .D (nx24133), .CLK (
        clk)) ;
    nand03 ix33152 (.Y (nx33151), .A0 (nx35181), .A1 (nx16674), .A2 (nx34815)) ;
    dff max_calc_reg_ans4_3 (.Q (max_calc_ans4_3), .QB (\$dummy [615]), .D (
        nx24123), .CLK (clk)) ;
    dff max_calc_reg_comparator_second_inp1_3 (.Q (
        max_calc_comparator_second_inp1_3), .QB (nx33160), .D (nx24153), .CLK (
        clk)) ;
    oai21 ix24154 (.Y (nx24153), .A0 (nx33160), .A1 (nx34815), .B0 (nx33163)) ;
    nand03 ix33164 (.Y (nx33163), .A0 (nx35181), .A1 (nx16710), .A2 (nx34815)) ;
    dff max_calc_reg_ans3_3 (.Q (max_calc_ans3_3), .QB (\$dummy [616]), .D (
        nx24143), .CLK (clk)) ;
    aoi22 ix33173 (.Y (nx33172), .A0 (nx33174), .A1 (
          max_calc_comparator_second_inp1_2), .B0 (nx16796), .B1 (nx16958)) ;
    dff max_calc_reg_comparator_second_inp2_2 (.Q (\$dummy [617]), .QB (nx33174)
        , .D (nx24173), .CLK (clk)) ;
    oai21 ix24174 (.Y (nx24173), .A0 (nx33174), .A1 (nx34815), .B0 (nx33177)) ;
    nand03 ix33178 (.Y (nx33177), .A0 (nx35181), .A1 (nx16748), .A2 (nx34817)) ;
    dff max_calc_reg_ans4_2 (.Q (max_calc_ans4_2), .QB (nx33184), .D (nx24163), 
        .CLK (clk)) ;
    oai21 ix24194 (.Y (nx24193), .A0 (nx33188), .A1 (nx34817), .B0 (nx33190)) ;
    dff max_calc_reg_comparator_second_inp1_2 (.Q (
        max_calc_comparator_second_inp1_2), .QB (nx33188), .D (nx24193), .CLK (
        clk)) ;
    nand03 ix33191 (.Y (nx33190), .A0 (nx35181), .A1 (nx16784), .A2 (nx34817)) ;
    dff max_calc_reg_ans3_2 (.Q (max_calc_ans3_2), .QB (nx33197), .D (nx24183), 
        .CLK (clk)) ;
    oai21 ix16959 (.Y (nx16958), .A0 (max_calc_comparator_second_inp2_1), .A1 (
          nx33214), .B0 (nx33226)) ;
    oai21 ix24214 (.Y (nx24213), .A0 (nx33203), .A1 (nx34817), .B0 (nx33205)) ;
    dff max_calc_reg_comparator_second_inp2_1 (.Q (
        max_calc_comparator_second_inp2_1), .QB (nx33203), .D (nx24213), .CLK (
        clk)) ;
    nand03 ix33206 (.Y (nx33205), .A0 (nx35181), .A1 (nx16822), .A2 (nx34817)) ;
    dff max_calc_reg_ans4_1 (.Q (max_calc_ans4_1), .QB (\$dummy [618]), .D (
        nx24203), .CLK (clk)) ;
    dff max_calc_reg_comparator_second_inp1_1 (.Q (\$dummy [619]), .QB (nx33214)
        , .D (nx24233), .CLK (clk)) ;
    oai21 ix24234 (.Y (nx24233), .A0 (nx33214), .A1 (nx34817), .B0 (nx33217)) ;
    nand03 ix33218 (.Y (nx33217), .A0 (nx35959), .A1 (nx16858), .A2 (nx34817)) ;
    dff max_calc_reg_ans3_1 (.Q (max_calc_ans3_1), .QB (\$dummy [620]), .D (
        nx24223), .CLK (clk)) ;
    oai21 ix33227 (.Y (nx33226), .A0 (nx30546), .A1 (
          max_calc_comparator_second_inp1_0), .B0 (nx16870)) ;
    oai21 ix24294 (.Y (nx24293), .A0 (nx33232), .A1 (nx34819), .B0 (nx33234)) ;
    dff max_calc_reg_comparator_second_inp2_15 (.Q (\$dummy [621]), .QB (nx33232
        ), .D (nx24293), .CLK (clk)) ;
    nand03 ix33235 (.Y (nx33234), .A0 (nx35959), .A1 (nx17088), .A2 (nx34819)) ;
    dffr labelsregfile_label4_loop1_15_fx_reg_q (.Q (label_4_output[15]), .QB (
         \$dummy [622]), .D (nx14963), .CLK (clk), .R (rst)) ;
    latch lat_label_4_input_15 (.Q (label_4_input_15), .D (nx2212), .CLK (
          nx34547)) ;
    dffr reg_label_4_input_state_machine_15 (.Q (label_4_input_state_machine_15)
         , .QB (\$dummy [623]), .D (nx14123), .CLK (clk), .R (rst)) ;
    xnor2 ix2209 (.Y (nx2208), .A0 (nx2204), .A1 (nx33246)) ;
    oai22 ix2205 (.Y (nx2204), .A0 (nx32486), .A1 (nx32658), .B0 (nx32660), .B1 (
          nx30968)) ;
    dff max_calc_reg_ans4_15 (.Q (max_calc_ans4_15), .QB (\$dummy [624]), .D (
        nx24283), .CLK (clk)) ;
    oai21 ix24314 (.Y (nx24313), .A0 (nx33257), .A1 (nx34819), .B0 (nx33259)) ;
    dff max_calc_reg_comparator_second_inp1_15 (.Q (\$dummy [625]), .QB (nx33257
        ), .D (nx24313), .CLK (clk)) ;
    nand03 ix33260 (.Y (nx33259), .A0 (nx35959), .A1 (nx17124), .A2 (nx34819)) ;
    dffr labelsregfile_label3_loop1_15_fx_reg_q (.Q (label_3_output[15]), .QB (
         \$dummy [626]), .D (nx15813), .CLK (clk), .R (rst)) ;
    latch lat_label_3_input_15 (.Q (label_3_input_15), .D (nx3550), .CLK (
          nx34547)) ;
    dffr reg_label_3_input_state_machine_15 (.Q (label_3_input_state_machine_15)
         , .QB (\$dummy [627]), .D (nx14973), .CLK (clk), .R (rst)) ;
    xnor2 ix3547 (.Y (nx3546), .A0 (nx3542), .A1 (nx33271)) ;
    oai22 ix3543 (.Y (nx3542), .A0 (nx32682), .A1 (nx32854), .B0 (nx32856), .B1 (
          nx29039)) ;
    dff max_calc_reg_ans3_15 (.Q (max_calc_ans3_15), .QB (\$dummy [628]), .D (
        nx24303), .CLK (clk)) ;
    dff max_calc_reg_ans7_0 (.Q (max_calc_ans7_0), .QB (\$dummy [629]), .D (
        nx25463), .CLK (clk)) ;
    dff max_calc_reg_ans8_0 (.Q (max_calc_ans8_0), .QB (\$dummy [630]), .D (
        nx25453), .CLK (clk)) ;
    xnor2 ix19143 (.Y (nx13373), .A0 (nx33290), .A1 (nx19140)) ;
    aoi22 ix33291 (.Y (nx33290), .A0 (nx33292), .A1 (
          max_calc_comparator_first_inp1_14), .B0 (nx17256), .B1 (nx19010)) ;
    dffr labelsregfile_label2_loop1_14_fx_reg_q (.Q (label_2_output[14]), .QB (
         nx33479), .D (nx16653), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_14 (.Q (label_2_input_14), .D (nx4862), .CLK (
          nx34551)) ;
    dffr reg_label_2_input_state_machine_14 (.Q (label_2_input_state_machine_14)
         , .QB (\$dummy [631]), .D (nx16643), .CLK (clk), .R (rst)) ;
    xor2 ix4859 (.Y (nx4858), .A0 (nx33305), .A1 (nx33477)) ;
    aoi22 ix33306 (.Y (nx33305), .A0 (label_2_output[13]), .A1 (
          booth_booth_integration_output_1_13), .B0 (nx4816), .B1 (nx13063)) ;
    dffr labelsregfile_label2_loop1_13_fx_reg_q (.Q (label_2_output[13]), .QB (
         \$dummy [632]), .D (nx16633), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_13 (.Q (label_2_input_13), .D (nx4830), .CLK (
          nx34551)) ;
    dffr reg_label_2_input_state_machine_13 (.Q (label_2_input_state_machine_13)
         , .QB (\$dummy [633]), .D (nx16623), .CLK (clk), .R (rst)) ;
    xnor2 ix4827 (.Y (nx4826), .A0 (nx4816), .A1 (nx33473)) ;
    oai22 ix4817 (.Y (nx4816), .A0 (nx33316), .A1 (nx33462), .B0 (nx33472), .B1 (
          nx28598)) ;
    aoi22 ix33317 (.Y (nx33316), .A0 (label_2_output[11]), .A1 (
          booth_booth_integration_output_1_11), .B0 (nx4752), .B1 (nx13059)) ;
    dffr labelsregfile_label2_loop1_11_fx_reg_q (.Q (label_2_output[11]), .QB (
         \$dummy [634]), .D (nx16593), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_11 (.Q (label_2_input_11), .D (nx4766), .CLK (
          nx34551)) ;
    dffr reg_label_2_input_state_machine_11 (.Q (label_2_input_state_machine_11)
         , .QB (\$dummy [635]), .D (nx16583), .CLK (clk), .R (rst)) ;
    xnor2 ix4763 (.Y (nx4762), .A0 (nx4752), .A1 (nx33458)) ;
    oai22 ix4753 (.Y (nx4752), .A0 (nx33327), .A1 (nx33447), .B0 (nx33457), .B1 (
          nx28600)) ;
    aoi22 ix33328 (.Y (nx33327), .A0 (label_2_output[9]), .A1 (
          booth_booth_integration_output_1_9), .B0 (nx4688), .B1 (nx13055)) ;
    dffr labelsregfile_label2_loop1_9_fx_reg_q (.Q (label_2_output[9]), .QB (
         \$dummy [636]), .D (nx16553), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_9 (.Q (label_2_input_9), .D (nx4702), .CLK (nx34549)
          ) ;
    dffr reg_label_2_input_state_machine_9 (.Q (label_2_input_state_machine_9), 
         .QB (\$dummy [637]), .D (nx16543), .CLK (clk), .R (rst)) ;
    xnor2 ix4699 (.Y (nx4698), .A0 (nx4688), .A1 (nx33443)) ;
    oai22 ix4689 (.Y (nx4688), .A0 (nx33338), .A1 (nx33432), .B0 (nx33442), .B1 (
          nx28602)) ;
    aoi22 ix33339 (.Y (nx33338), .A0 (label_2_output[7]), .A1 (
          booth_booth_integration_output_1_7), .B0 (nx4624), .B1 (nx13051)) ;
    dffr labelsregfile_label2_loop1_7_fx_reg_q (.Q (label_2_output[7]), .QB (
         \$dummy [638]), .D (nx16513), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_7 (.Q (label_2_input_7), .D (nx4638), .CLK (nx34549)
          ) ;
    dffr reg_label_2_input_state_machine_7 (.Q (label_2_input_state_machine_7), 
         .QB (\$dummy [639]), .D (nx16503), .CLK (clk), .R (rst)) ;
    xnor2 ix4635 (.Y (nx4634), .A0 (nx4624), .A1 (nx33428)) ;
    oai22 ix4625 (.Y (nx4624), .A0 (nx33349), .A1 (nx33417), .B0 (nx33427), .B1 (
          nx28604)) ;
    aoi22 ix33350 (.Y (nx33349), .A0 (label_2_output[5]), .A1 (
          booth_booth_integration_output_1_5), .B0 (nx4560), .B1 (nx13049)) ;
    dffr labelsregfile_label2_loop1_5_fx_reg_q (.Q (label_2_output[5]), .QB (
         \$dummy [640]), .D (nx16473), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_5 (.Q (label_2_input_5), .D (nx4574), .CLK (nx34549)
          ) ;
    dffr reg_label_2_input_state_machine_5 (.Q (label_2_input_state_machine_5), 
         .QB (\$dummy [641]), .D (nx16463), .CLK (clk), .R (rst)) ;
    xnor2 ix4571 (.Y (nx4570), .A0 (nx4560), .A1 (nx33413)) ;
    oai22 ix4561 (.Y (nx4560), .A0 (nx33360), .A1 (nx33402), .B0 (nx33412), .B1 (
          nx28606)) ;
    aoi22 ix33361 (.Y (nx33360), .A0 (label_2_output[3]), .A1 (
          booth_booth_integration_output_1_3), .B0 (nx4496), .B1 (nx13045)) ;
    dffr labelsregfile_label2_loop1_3_fx_reg_q (.Q (label_2_output[3]), .QB (
         \$dummy [642]), .D (nx16433), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_3 (.Q (label_2_input_3), .D (nx4510), .CLK (nx34547)
          ) ;
    dffr reg_label_2_input_state_machine_3 (.Q (label_2_input_state_machine_3), 
         .QB (\$dummy [643]), .D (nx16423), .CLK (clk), .R (rst)) ;
    xnor2 ix4507 (.Y (nx4506), .A0 (nx4496), .A1 (nx33398)) ;
    oai22 ix4497 (.Y (nx4496), .A0 (nx33371), .A1 (nx33387), .B0 (nx33397), .B1 (
          nx28608)) ;
    aoi32 ix33372 (.Y (nx33371), .A0 (label_2_output[0]), .A1 (nx35727), .A2 (
          nx13042), .B0 (label_2_output[1]), .B1 (
          booth_booth_integration_output_1_1)) ;
    dffr labelsregfile_label2_loop1_1_fx_reg_q (.Q (label_2_output[1]), .QB (
         \$dummy [644]), .D (nx16393), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_1 (.Q (label_2_input_1), .D (nx4446), .CLK (nx34547)
          ) ;
    dffr reg_label_2_input_state_machine_1 (.Q (label_2_input_state_machine_1), 
         .QB (\$dummy [645]), .D (nx16383), .CLK (clk), .R (rst)) ;
    xor2 ix4443 (.Y (nx4442), .A0 (nx33382), .A1 (nx33384)) ;
    nand02 ix33383 (.Y (nx33382), .A0 (label_2_output[0]), .A1 (nx35727)) ;
    xnor2 ix33385 (.Y (nx33384), .A0 (booth_booth_integration_output_1_1), .A1 (
          label_2_output[1])) ;
    dffr labelsregfile_label2_loop1_2_fx_reg_q (.Q (label_2_output[2]), .QB (
         nx33397), .D (nx16413), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_2 (.Q (label_2_input_2), .D (nx4478), .CLK (nx34547)
          ) ;
    dffr reg_label_2_input_state_machine_2 (.Q (label_2_input_state_machine_2), 
         .QB (\$dummy [646]), .D (nx16403), .CLK (clk), .R (rst)) ;
    xor2 ix4475 (.Y (nx4474), .A0 (nx33371), .A1 (nx33387)) ;
    xnor2 ix33399 (.Y (nx33398), .A0 (booth_booth_integration_output_1_3), .A1 (
          label_2_output[3])) ;
    dffr labelsregfile_label2_loop1_4_fx_reg_q (.Q (label_2_output[4]), .QB (
         nx33412), .D (nx16453), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_4 (.Q (label_2_input_4), .D (nx4542), .CLK (nx34549)
          ) ;
    dffr reg_label_2_input_state_machine_4 (.Q (label_2_input_state_machine_4), 
         .QB (\$dummy [647]), .D (nx16443), .CLK (clk), .R (rst)) ;
    xor2 ix4539 (.Y (nx4538), .A0 (nx33360), .A1 (nx33402)) ;
    xnor2 ix33414 (.Y (nx33413), .A0 (booth_booth_integration_output_1_5), .A1 (
          label_2_output[5])) ;
    dffr labelsregfile_label2_loop1_6_fx_reg_q (.Q (label_2_output[6]), .QB (
         nx33427), .D (nx16493), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_6 (.Q (label_2_input_6), .D (nx4606), .CLK (nx34549)
          ) ;
    dffr reg_label_2_input_state_machine_6 (.Q (label_2_input_state_machine_6), 
         .QB (\$dummy [648]), .D (nx16483), .CLK (clk), .R (rst)) ;
    xor2 ix4603 (.Y (nx4602), .A0 (nx33349), .A1 (nx33417)) ;
    xnor2 ix33429 (.Y (nx33428), .A0 (booth_booth_integration_output_1_7), .A1 (
          label_2_output[7])) ;
    dffr labelsregfile_label2_loop1_8_fx_reg_q (.Q (label_2_output[8]), .QB (
         nx33442), .D (nx16533), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_8 (.Q (label_2_input_8), .D (nx4670), .CLK (nx34549)
          ) ;
    dffr reg_label_2_input_state_machine_8 (.Q (label_2_input_state_machine_8), 
         .QB (\$dummy [649]), .D (nx16523), .CLK (clk), .R (rst)) ;
    xor2 ix4667 (.Y (nx4666), .A0 (nx33338), .A1 (nx33432)) ;
    xnor2 ix33444 (.Y (nx33443), .A0 (booth_booth_integration_output_1_9), .A1 (
          label_2_output[9])) ;
    dffr labelsregfile_label2_loop1_10_fx_reg_q (.Q (label_2_output[10]), .QB (
         nx33457), .D (nx16573), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_10 (.Q (label_2_input_10), .D (nx4734), .CLK (
          nx34549)) ;
    dffr reg_label_2_input_state_machine_10 (.Q (label_2_input_state_machine_10)
         , .QB (\$dummy [650]), .D (nx16563), .CLK (clk), .R (rst)) ;
    xor2 ix4731 (.Y (nx4730), .A0 (nx33327), .A1 (nx33447)) ;
    xnor2 ix33459 (.Y (nx33458), .A0 (booth_booth_integration_output_1_11), .A1 (
          label_2_output[11])) ;
    dffr labelsregfile_label2_loop1_12_fx_reg_q (.Q (label_2_output[12]), .QB (
         nx33472), .D (nx16613), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_12 (.Q (label_2_input_12), .D (nx4798), .CLK (
          nx34551)) ;
    dffr reg_label_2_input_state_machine_12 (.Q (label_2_input_state_machine_12)
         , .QB (\$dummy [651]), .D (nx16603), .CLK (clk), .R (rst)) ;
    xor2 ix4795 (.Y (nx4794), .A0 (nx33316), .A1 (nx33462)) ;
    xnor2 ix33474 (.Y (nx33473), .A0 (booth_booth_integration_output_1_13), .A1 (
          label_2_output[13])) ;
    dff max_calc_reg_ans2_14 (.Q (max_calc_ans2_14), .QB (\$dummy [652]), .D (
        nx24323), .CLK (clk)) ;
    dff max_calc_reg_ans7_14 (.Q (max_calc_ans7_14), .QB (\$dummy [653]), .D (
        nx24383), .CLK (clk)) ;
    dff max_calc_reg_ans8_14 (.Q (max_calc_ans8_14), .QB (\$dummy [654]), .D (
        nx24373), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_14 (.Q (
        max_calc_comparator_first_inp1_14), .QB (\$dummy [655]), .D (nx24363), .CLK (
        clk)) ;
    dffr labelsregfile_label1_loop1_14_fx_reg_q (.Q (label_1_output[14]), .QB (
         nx33677), .D (nx17503), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_14 (.Q (label_1_input_14), .D (nx6200), .CLK (
          nx34555)) ;
    dffr reg_label_1_input_state_machine_14 (.Q (label_1_input_state_machine_14)
         , .QB (\$dummy [656]), .D (nx17493), .CLK (clk), .R (rst)) ;
    xor2 ix6197 (.Y (nx6196), .A0 (nx33503), .A1 (nx33675)) ;
    aoi22 ix33504 (.Y (nx33503), .A0 (label_1_output[13]), .A1 (
          booth_booth_integration_output_0_13), .B0 (nx6154), .B1 (nx13114)) ;
    dffr labelsregfile_label1_loop1_13_fx_reg_q (.Q (label_1_output[13]), .QB (
         \$dummy [657]), .D (nx17483), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_13 (.Q (label_1_input_13), .D (nx6168), .CLK (
          nx34555)) ;
    dffr reg_label_1_input_state_machine_13 (.Q (label_1_input_state_machine_13)
         , .QB (\$dummy [658]), .D (nx17473), .CLK (clk), .R (rst)) ;
    xnor2 ix6165 (.Y (nx6164), .A0 (nx6154), .A1 (nx33671)) ;
    oai22 ix6155 (.Y (nx6154), .A0 (nx33514), .A1 (nx33660), .B0 (nx33670), .B1 (
          nx26638)) ;
    aoi22 ix33515 (.Y (nx33514), .A0 (label_1_output[11]), .A1 (
          booth_booth_integration_output_0_11), .B0 (nx6090), .B1 (nx13111)) ;
    dffr labelsregfile_label1_loop1_11_fx_reg_q (.Q (label_1_output[11]), .QB (
         \$dummy [659]), .D (nx17443), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_11 (.Q (label_1_input_11), .D (nx6104), .CLK (
          nx34555)) ;
    dffr reg_label_1_input_state_machine_11 (.Q (label_1_input_state_machine_11)
         , .QB (\$dummy [660]), .D (nx17433), .CLK (clk), .R (rst)) ;
    xnor2 ix6101 (.Y (nx6100), .A0 (nx6090), .A1 (nx33656)) ;
    oai22 ix6091 (.Y (nx6090), .A0 (nx33525), .A1 (nx33645), .B0 (nx33655), .B1 (
          nx26640)) ;
    aoi22 ix33526 (.Y (nx33525), .A0 (label_1_output[9]), .A1 (
          booth_booth_integration_output_0_9), .B0 (nx6026), .B1 (nx13107)) ;
    dffr labelsregfile_label1_loop1_9_fx_reg_q (.Q (label_1_output[9]), .QB (
         \$dummy [661]), .D (nx17403), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_9 (.Q (label_1_input_9), .D (nx6040), .CLK (nx34553)
          ) ;
    dffr reg_label_1_input_state_machine_9 (.Q (label_1_input_state_machine_9), 
         .QB (\$dummy [662]), .D (nx17393), .CLK (clk), .R (rst)) ;
    xnor2 ix6037 (.Y (nx6036), .A0 (nx6026), .A1 (nx33641)) ;
    oai22 ix6027 (.Y (nx6026), .A0 (nx33536), .A1 (nx33630), .B0 (nx33640), .B1 (
          nx26642)) ;
    aoi22 ix33537 (.Y (nx33536), .A0 (label_1_output[7]), .A1 (
          booth_booth_integration_output_0_7), .B0 (nx5962), .B1 (nx13103)) ;
    dffr labelsregfile_label1_loop1_7_fx_reg_q (.Q (label_1_output[7]), .QB (
         \$dummy [663]), .D (nx17363), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_7 (.Q (label_1_input_7), .D (nx5976), .CLK (nx34553)
          ) ;
    dffr reg_label_1_input_state_machine_7 (.Q (label_1_input_state_machine_7), 
         .QB (\$dummy [664]), .D (nx17353), .CLK (clk), .R (rst)) ;
    xnor2 ix5973 (.Y (nx5972), .A0 (nx5962), .A1 (nx33626)) ;
    oai22 ix5963 (.Y (nx5962), .A0 (nx33547), .A1 (nx33615), .B0 (nx33625), .B1 (
          nx26644)) ;
    aoi22 ix33548 (.Y (nx33547), .A0 (label_1_output[5]), .A1 (
          booth_booth_integration_output_0_5), .B0 (nx5898), .B1 (nx13099)) ;
    dffr labelsregfile_label1_loop1_5_fx_reg_q (.Q (label_1_output[5]), .QB (
         \$dummy [665]), .D (nx17323), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_5 (.Q (label_1_input_5), .D (nx5912), .CLK (nx34553)
          ) ;
    dffr reg_label_1_input_state_machine_5 (.Q (label_1_input_state_machine_5), 
         .QB (\$dummy [666]), .D (nx17313), .CLK (clk), .R (rst)) ;
    xnor2 ix5909 (.Y (nx5908), .A0 (nx5898), .A1 (nx33611)) ;
    oai22 ix5899 (.Y (nx5898), .A0 (nx33558), .A1 (nx33600), .B0 (nx33610), .B1 (
          nx26646)) ;
    aoi22 ix33559 (.Y (nx33558), .A0 (label_1_output[3]), .A1 (
          booth_booth_integration_output_0_3), .B0 (nx5834), .B1 (nx13097)) ;
    dffr labelsregfile_label1_loop1_3_fx_reg_q (.Q (label_1_output[3]), .QB (
         \$dummy [667]), .D (nx17283), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_3 (.Q (label_1_input_3), .D (nx5848), .CLK (nx34551)
          ) ;
    dffr reg_label_1_input_state_machine_3 (.Q (label_1_input_state_machine_3), 
         .QB (\$dummy [668]), .D (nx17273), .CLK (clk), .R (rst)) ;
    xnor2 ix5845 (.Y (nx5844), .A0 (nx5834), .A1 (nx33596)) ;
    oai22 ix5835 (.Y (nx5834), .A0 (nx33569), .A1 (nx33585), .B0 (nx33595), .B1 (
          nx26648)) ;
    aoi32 ix33570 (.Y (nx33569), .A0 (label_1_output[0]), .A1 (nx35731), .A2 (
          nx13093), .B0 (label_1_output[1]), .B1 (
          booth_booth_integration_output_0_1)) ;
    dffr labelsregfile_label1_loop1_1_fx_reg_q (.Q (label_1_output[1]), .QB (
         \$dummy [669]), .D (nx17243), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_1 (.Q (label_1_input_1), .D (nx5784), .CLK (nx34551)
          ) ;
    dffr reg_label_1_input_state_machine_1 (.Q (label_1_input_state_machine_1), 
         .QB (\$dummy [670]), .D (nx17233), .CLK (clk), .R (rst)) ;
    xor2 ix5781 (.Y (nx5780), .A0 (nx33580), .A1 (nx33582)) ;
    nand02 ix33581 (.Y (nx33580), .A0 (label_1_output[0]), .A1 (nx35731)) ;
    xnor2 ix33583 (.Y (nx33582), .A0 (booth_booth_integration_output_0_1), .A1 (
          label_1_output[1])) ;
    dffr labelsregfile_label1_loop1_2_fx_reg_q (.Q (label_1_output[2]), .QB (
         nx33595), .D (nx17263), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_2 (.Q (label_1_input_2), .D (nx5816), .CLK (nx34551)
          ) ;
    dffr reg_label_1_input_state_machine_2 (.Q (label_1_input_state_machine_2), 
         .QB (\$dummy [671]), .D (nx17253), .CLK (clk), .R (rst)) ;
    xor2 ix5813 (.Y (nx5812), .A0 (nx33569), .A1 (nx33585)) ;
    xnor2 ix33597 (.Y (nx33596), .A0 (booth_booth_integration_output_0_3), .A1 (
          label_1_output[3])) ;
    dffr labelsregfile_label1_loop1_4_fx_reg_q (.Q (label_1_output[4]), .QB (
         nx33610), .D (nx17303), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_4 (.Q (label_1_input_4), .D (nx5880), .CLK (nx34553)
          ) ;
    dffr reg_label_1_input_state_machine_4 (.Q (label_1_input_state_machine_4), 
         .QB (\$dummy [672]), .D (nx17293), .CLK (clk), .R (rst)) ;
    xor2 ix5877 (.Y (nx5876), .A0 (nx33558), .A1 (nx33600)) ;
    xnor2 ix33612 (.Y (nx33611), .A0 (booth_booth_integration_output_0_5), .A1 (
          label_1_output[5])) ;
    dffr labelsregfile_label1_loop1_6_fx_reg_q (.Q (label_1_output[6]), .QB (
         nx33625), .D (nx17343), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_6 (.Q (label_1_input_6), .D (nx5944), .CLK (nx34553)
          ) ;
    dffr reg_label_1_input_state_machine_6 (.Q (label_1_input_state_machine_6), 
         .QB (\$dummy [673]), .D (nx17333), .CLK (clk), .R (rst)) ;
    xor2 ix5941 (.Y (nx5940), .A0 (nx33547), .A1 (nx33615)) ;
    xnor2 ix33627 (.Y (nx33626), .A0 (booth_booth_integration_output_0_7), .A1 (
          label_1_output[7])) ;
    dffr labelsregfile_label1_loop1_8_fx_reg_q (.Q (label_1_output[8]), .QB (
         nx33640), .D (nx17383), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_8 (.Q (label_1_input_8), .D (nx6008), .CLK (nx34553)
          ) ;
    dffr reg_label_1_input_state_machine_8 (.Q (label_1_input_state_machine_8), 
         .QB (\$dummy [674]), .D (nx17373), .CLK (clk), .R (rst)) ;
    xor2 ix6005 (.Y (nx6004), .A0 (nx33536), .A1 (nx33630)) ;
    xnor2 ix33642 (.Y (nx33641), .A0 (booth_booth_integration_output_0_9), .A1 (
          label_1_output[9])) ;
    dffr labelsregfile_label1_loop1_10_fx_reg_q (.Q (label_1_output[10]), .QB (
         nx33655), .D (nx17423), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_10 (.Q (label_1_input_10), .D (nx6072), .CLK (
          nx34553)) ;
    dffr reg_label_1_input_state_machine_10 (.Q (label_1_input_state_machine_10)
         , .QB (\$dummy [675]), .D (nx17413), .CLK (clk), .R (rst)) ;
    xor2 ix6069 (.Y (nx6068), .A0 (nx33525), .A1 (nx33645)) ;
    xnor2 ix33657 (.Y (nx33656), .A0 (booth_booth_integration_output_0_11), .A1 (
          label_1_output[11])) ;
    dffr labelsregfile_label1_loop1_12_fx_reg_q (.Q (label_1_output[12]), .QB (
         nx33670), .D (nx17463), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_12 (.Q (label_1_input_12), .D (nx6136), .CLK (
          nx34555)) ;
    dffr reg_label_1_input_state_machine_12 (.Q (label_1_input_state_machine_12)
         , .QB (\$dummy [676]), .D (nx17453), .CLK (clk), .R (rst)) ;
    xor2 ix6133 (.Y (nx6132), .A0 (nx33514), .A1 (nx33660)) ;
    xnor2 ix33672 (.Y (nx33671), .A0 (booth_booth_integration_output_0_13), .A1 (
          label_1_output[13])) ;
    dff max_calc_reg_ans1_14 (.Q (max_calc_ans1_14), .QB (\$dummy [677]), .D (
        nx24333), .CLK (clk)) ;
    dff max_calc_reg_ans6_14 (.Q (max_calc_ans6_14), .QB (\$dummy [678]), .D (
        nx24343), .CLK (clk)) ;
    dff max_calc_reg_ans5_14 (.Q (max_calc_ans5_14), .QB (\$dummy [679]), .D (
        nx24353), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp2_14 (.Q (
        max_calc_comparator_first_inp2_14), .QB (nx33292), .D (nx24393), .CLK (
        clk)) ;
    oai22 ix19011 (.Y (nx19010), .A0 (nx33694), .A1 (nx33729), .B0 (
          max_calc_comparator_first_inp2_13), .B1 (nx33726)) ;
    dff max_calc_reg_comparator_first_inp2_13 (.Q (
        max_calc_comparator_first_inp2_13), .QB (\$dummy [680]), .D (nx24473), .CLK (
        clk)) ;
    dff max_calc_reg_ans2_13 (.Q (max_calc_ans2_13), .QB (\$dummy [681]), .D (
        nx24403), .CLK (clk)) ;
    dff max_calc_reg_ans7_13 (.Q (max_calc_ans7_13), .QB (\$dummy [682]), .D (
        nx24463), .CLK (clk)) ;
    dff max_calc_reg_ans8_13 (.Q (max_calc_ans8_13), .QB (\$dummy [683]), .D (
        nx24453), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_13 (.Q (
        max_calc_comparator_first_inp1_13), .QB (nx33726), .D (nx24443), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_13 (.Q (max_calc_ans1_13), .QB (\$dummy [684]), .D (
        nx24413), .CLK (clk)) ;
    dff max_calc_reg_ans6_13 (.Q (max_calc_ans6_13), .QB (\$dummy [685]), .D (
        nx24423), .CLK (clk)) ;
    dff max_calc_reg_ans5_13 (.Q (max_calc_ans5_13), .QB (\$dummy [686]), .D (
        nx24433), .CLK (clk)) ;
    aoi22 ix33730 (.Y (nx33729), .A0 (nx33731), .A1 (
          max_calc_comparator_first_inp1_12), .B0 (nx17500), .B1 (nx18994)) ;
    dff max_calc_reg_ans2_12 (.Q (max_calc_ans2_12), .QB (\$dummy [687]), .D (
        nx24483), .CLK (clk)) ;
    dff max_calc_reg_ans7_12 (.Q (max_calc_ans7_12), .QB (\$dummy [688]), .D (
        nx24543), .CLK (clk)) ;
    dff max_calc_reg_ans8_12 (.Q (max_calc_ans8_12), .QB (\$dummy [689]), .D (
        nx24533), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_12 (.Q (
        max_calc_comparator_first_inp1_12), .QB (\$dummy [690]), .D (nx24523), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_12 (.Q (max_calc_ans1_12), .QB (\$dummy [691]), .D (
        nx24493), .CLK (clk)) ;
    dff max_calc_reg_ans6_12 (.Q (max_calc_ans6_12), .QB (\$dummy [692]), .D (
        nx24503), .CLK (clk)) ;
    dff max_calc_reg_ans5_12 (.Q (max_calc_ans5_12), .QB (\$dummy [693]), .D (
        nx24513), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp2_12 (.Q (
        max_calc_comparator_first_inp2_12), .QB (nx33731), .D (nx24553), .CLK (
        clk)) ;
    oai22 ix18995 (.Y (nx18994), .A0 (nx33767), .A1 (nx33802), .B0 (
          max_calc_comparator_first_inp2_11), .B1 (nx33799)) ;
    dff max_calc_reg_comparator_first_inp2_11 (.Q (
        max_calc_comparator_first_inp2_11), .QB (\$dummy [694]), .D (nx24633), .CLK (
        clk)) ;
    dff max_calc_reg_ans2_11 (.Q (max_calc_ans2_11), .QB (\$dummy [695]), .D (
        nx24563), .CLK (clk)) ;
    dff max_calc_reg_ans7_11 (.Q (max_calc_ans7_11), .QB (\$dummy [696]), .D (
        nx24623), .CLK (clk)) ;
    dff max_calc_reg_ans8_11 (.Q (max_calc_ans8_11), .QB (\$dummy [697]), .D (
        nx24613), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_11 (.Q (
        max_calc_comparator_first_inp1_11), .QB (nx33799), .D (nx24603), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_11 (.Q (max_calc_ans1_11), .QB (\$dummy [698]), .D (
        nx24573), .CLK (clk)) ;
    dff max_calc_reg_ans6_11 (.Q (max_calc_ans6_11), .QB (\$dummy [699]), .D (
        nx24583), .CLK (clk)) ;
    dff max_calc_reg_ans5_11 (.Q (max_calc_ans5_11), .QB (\$dummy [700]), .D (
        nx24593), .CLK (clk)) ;
    aoi22 ix33803 (.Y (nx33802), .A0 (nx33804), .A1 (
          max_calc_comparator_first_inp1_10), .B0 (nx17744), .B1 (nx18978)) ;
    dff max_calc_reg_ans2_10 (.Q (max_calc_ans2_10), .QB (\$dummy [701]), .D (
        nx24643), .CLK (clk)) ;
    dff max_calc_reg_ans7_10 (.Q (max_calc_ans7_10), .QB (\$dummy [702]), .D (
        nx24703), .CLK (clk)) ;
    dff max_calc_reg_ans8_10 (.Q (max_calc_ans8_10), .QB (\$dummy [703]), .D (
        nx24693), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_10 (.Q (
        max_calc_comparator_first_inp1_10), .QB (\$dummy [704]), .D (nx24683), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_10 (.Q (max_calc_ans1_10), .QB (\$dummy [705]), .D (
        nx24653), .CLK (clk)) ;
    dff max_calc_reg_ans6_10 (.Q (max_calc_ans6_10), .QB (\$dummy [706]), .D (
        nx24663), .CLK (clk)) ;
    dff max_calc_reg_ans5_10 (.Q (max_calc_ans5_10), .QB (\$dummy [707]), .D (
        nx24673), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp2_10 (.Q (
        max_calc_comparator_first_inp2_10), .QB (nx33804), .D (nx24713), .CLK (
        clk)) ;
    oai22 ix18979 (.Y (nx18978), .A0 (nx33840), .A1 (nx33875), .B0 (
          max_calc_comparator_first_inp2_9), .B1 (nx33872)) ;
    dff max_calc_reg_comparator_first_inp2_9 (.Q (
        max_calc_comparator_first_inp2_9), .QB (\$dummy [708]), .D (nx24793), .CLK (
        clk)) ;
    dff max_calc_reg_ans2_9 (.Q (max_calc_ans2_9), .QB (\$dummy [709]), .D (
        nx24723), .CLK (clk)) ;
    dff max_calc_reg_ans7_9 (.Q (max_calc_ans7_9), .QB (\$dummy [710]), .D (
        nx24783), .CLK (clk)) ;
    dff max_calc_reg_ans8_9 (.Q (max_calc_ans8_9), .QB (\$dummy [711]), .D (
        nx24773), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_9 (.Q (
        max_calc_comparator_first_inp1_9), .QB (nx33872), .D (nx24763), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_9 (.Q (max_calc_ans1_9), .QB (\$dummy [712]), .D (
        nx24733), .CLK (clk)) ;
    dff max_calc_reg_ans6_9 (.Q (max_calc_ans6_9), .QB (\$dummy [713]), .D (
        nx24743), .CLK (clk)) ;
    dff max_calc_reg_ans5_9 (.Q (max_calc_ans5_9), .QB (\$dummy [714]), .D (
        nx24753), .CLK (clk)) ;
    aoi22 ix33876 (.Y (nx33875), .A0 (nx33877), .A1 (
          max_calc_comparator_first_inp1_8), .B0 (nx17988), .B1 (nx18962)) ;
    dff max_calc_reg_ans2_8 (.Q (max_calc_ans2_8), .QB (\$dummy [715]), .D (
        nx24803), .CLK (clk)) ;
    dff max_calc_reg_ans7_8 (.Q (max_calc_ans7_8), .QB (\$dummy [716]), .D (
        nx24863), .CLK (clk)) ;
    dff max_calc_reg_ans8_8 (.Q (max_calc_ans8_8), .QB (\$dummy [717]), .D (
        nx24853), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_8 (.Q (
        max_calc_comparator_first_inp1_8), .QB (\$dummy [718]), .D (nx24843), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_8 (.Q (max_calc_ans1_8), .QB (\$dummy [719]), .D (
        nx24813), .CLK (clk)) ;
    dff max_calc_reg_ans6_8 (.Q (max_calc_ans6_8), .QB (\$dummy [720]), .D (
        nx24823), .CLK (clk)) ;
    dff max_calc_reg_ans5_8 (.Q (max_calc_ans5_8), .QB (\$dummy [721]), .D (
        nx24833), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp2_8 (.Q (
        max_calc_comparator_first_inp2_8), .QB (nx33877), .D (nx24873), .CLK (
        clk)) ;
    oai22 ix18963 (.Y (nx18962), .A0 (nx33913), .A1 (nx33948), .B0 (
          max_calc_comparator_first_inp2_7), .B1 (nx33945)) ;
    dff max_calc_reg_comparator_first_inp2_7 (.Q (
        max_calc_comparator_first_inp2_7), .QB (\$dummy [722]), .D (nx24953), .CLK (
        clk)) ;
    dff max_calc_reg_ans2_7 (.Q (max_calc_ans2_7), .QB (\$dummy [723]), .D (
        nx24883), .CLK (clk)) ;
    dff max_calc_reg_ans7_7 (.Q (max_calc_ans7_7), .QB (\$dummy [724]), .D (
        nx24943), .CLK (clk)) ;
    dff max_calc_reg_ans8_7 (.Q (max_calc_ans8_7), .QB (\$dummy [725]), .D (
        nx24933), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_7 (.Q (
        max_calc_comparator_first_inp1_7), .QB (nx33945), .D (nx24923), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_7 (.Q (max_calc_ans1_7), .QB (\$dummy [726]), .D (
        nx24893), .CLK (clk)) ;
    dff max_calc_reg_ans6_7 (.Q (max_calc_ans6_7), .QB (\$dummy [727]), .D (
        nx24903), .CLK (clk)) ;
    dff max_calc_reg_ans5_7 (.Q (max_calc_ans5_7), .QB (\$dummy [728]), .D (
        nx24913), .CLK (clk)) ;
    aoi22 ix33949 (.Y (nx33948), .A0 (nx33950), .A1 (
          max_calc_comparator_first_inp1_6), .B0 (nx18232), .B1 (nx18946)) ;
    dff max_calc_reg_ans2_6 (.Q (max_calc_ans2_6), .QB (\$dummy [729]), .D (
        nx24963), .CLK (clk)) ;
    dff max_calc_reg_ans7_6 (.Q (max_calc_ans7_6), .QB (\$dummy [730]), .D (
        nx25023), .CLK (clk)) ;
    dff max_calc_reg_ans8_6 (.Q (max_calc_ans8_6), .QB (\$dummy [731]), .D (
        nx25013), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_6 (.Q (
        max_calc_comparator_first_inp1_6), .QB (\$dummy [732]), .D (nx25003), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_6 (.Q (max_calc_ans1_6), .QB (\$dummy [733]), .D (
        nx24973), .CLK (clk)) ;
    dff max_calc_reg_ans6_6 (.Q (max_calc_ans6_6), .QB (\$dummy [734]), .D (
        nx24983), .CLK (clk)) ;
    dff max_calc_reg_ans5_6 (.Q (max_calc_ans5_6), .QB (\$dummy [735]), .D (
        nx24993), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp2_6 (.Q (
        max_calc_comparator_first_inp2_6), .QB (nx33950), .D (nx25033), .CLK (
        clk)) ;
    oai22 ix18947 (.Y (nx18946), .A0 (nx33986), .A1 (nx34021), .B0 (
          max_calc_comparator_first_inp2_5), .B1 (nx34018)) ;
    dff max_calc_reg_comparator_first_inp2_5 (.Q (
        max_calc_comparator_first_inp2_5), .QB (\$dummy [736]), .D (nx25113), .CLK (
        clk)) ;
    dff max_calc_reg_ans2_5 (.Q (max_calc_ans2_5), .QB (\$dummy [737]), .D (
        nx25043), .CLK (clk)) ;
    dff max_calc_reg_ans7_5 (.Q (max_calc_ans7_5), .QB (\$dummy [738]), .D (
        nx25103), .CLK (clk)) ;
    dff max_calc_reg_ans8_5 (.Q (max_calc_ans8_5), .QB (\$dummy [739]), .D (
        nx25093), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_5 (.Q (
        max_calc_comparator_first_inp1_5), .QB (nx34018), .D (nx25083), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_5 (.Q (max_calc_ans1_5), .QB (\$dummy [740]), .D (
        nx25053), .CLK (clk)) ;
    dff max_calc_reg_ans6_5 (.Q (max_calc_ans6_5), .QB (\$dummy [741]), .D (
        nx25063), .CLK (clk)) ;
    dff max_calc_reg_ans5_5 (.Q (max_calc_ans5_5), .QB (\$dummy [742]), .D (
        nx25073), .CLK (clk)) ;
    aoi22 ix34022 (.Y (nx34021), .A0 (nx34023), .A1 (
          max_calc_comparator_first_inp1_4), .B0 (nx18476), .B1 (nx18930)) ;
    dff max_calc_reg_ans2_4 (.Q (max_calc_ans2_4), .QB (\$dummy [743]), .D (
        nx25123), .CLK (clk)) ;
    dff max_calc_reg_ans7_4 (.Q (max_calc_ans7_4), .QB (\$dummy [744]), .D (
        nx25183), .CLK (clk)) ;
    dff max_calc_reg_ans8_4 (.Q (max_calc_ans8_4), .QB (\$dummy [745]), .D (
        nx25173), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_4 (.Q (
        max_calc_comparator_first_inp1_4), .QB (\$dummy [746]), .D (nx25163), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_4 (.Q (max_calc_ans1_4), .QB (\$dummy [747]), .D (
        nx25133), .CLK (clk)) ;
    dff max_calc_reg_ans6_4 (.Q (max_calc_ans6_4), .QB (\$dummy [748]), .D (
        nx25143), .CLK (clk)) ;
    dff max_calc_reg_ans5_4 (.Q (max_calc_ans5_4), .QB (\$dummy [749]), .D (
        nx25153), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp2_4 (.Q (
        max_calc_comparator_first_inp2_4), .QB (nx34023), .D (nx25193), .CLK (
        clk)) ;
    oai22 ix18931 (.Y (nx18930), .A0 (nx34059), .A1 (nx34094), .B0 (
          max_calc_comparator_first_inp2_3), .B1 (nx34091)) ;
    dff max_calc_reg_comparator_first_inp2_3 (.Q (
        max_calc_comparator_first_inp2_3), .QB (\$dummy [750]), .D (nx25273), .CLK (
        clk)) ;
    dff max_calc_reg_ans2_3 (.Q (max_calc_ans2_3), .QB (\$dummy [751]), .D (
        nx25203), .CLK (clk)) ;
    dff max_calc_reg_ans7_3 (.Q (max_calc_ans7_3), .QB (\$dummy [752]), .D (
        nx25263), .CLK (clk)) ;
    dff max_calc_reg_ans8_3 (.Q (max_calc_ans8_3), .QB (\$dummy [753]), .D (
        nx25253), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_3 (.Q (
        max_calc_comparator_first_inp1_3), .QB (nx34091), .D (nx25243), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_3 (.Q (max_calc_ans1_3), .QB (\$dummy [754]), .D (
        nx25213), .CLK (clk)) ;
    dff max_calc_reg_ans6_3 (.Q (max_calc_ans6_3), .QB (\$dummy [755]), .D (
        nx25223), .CLK (clk)) ;
    dff max_calc_reg_ans5_3 (.Q (max_calc_ans5_3), .QB (\$dummy [756]), .D (
        nx25233), .CLK (clk)) ;
    aoi22 ix34095 (.Y (nx34094), .A0 (nx34096), .A1 (
          max_calc_comparator_first_inp1_2), .B0 (nx18720), .B1 (nx18914)) ;
    dff max_calc_reg_ans2_2 (.Q (max_calc_ans2_2), .QB (\$dummy [757]), .D (
        nx25283), .CLK (clk)) ;
    dff max_calc_reg_ans7_2 (.Q (max_calc_ans7_2), .QB (\$dummy [758]), .D (
        nx25343), .CLK (clk)) ;
    dff max_calc_reg_ans8_2 (.Q (max_calc_ans8_2), .QB (\$dummy [759]), .D (
        nx25333), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_2 (.Q (
        max_calc_comparator_first_inp1_2), .QB (\$dummy [760]), .D (nx25323), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_2 (.Q (max_calc_ans1_2), .QB (\$dummy [761]), .D (
        nx25293), .CLK (clk)) ;
    dff max_calc_reg_ans6_2 (.Q (max_calc_ans6_2), .QB (\$dummy [762]), .D (
        nx25303), .CLK (clk)) ;
    dff max_calc_reg_ans5_2 (.Q (max_calc_ans5_2), .QB (\$dummy [763]), .D (
        nx25313), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp2_2 (.Q (
        max_calc_comparator_first_inp2_2), .QB (nx34096), .D (nx25353), .CLK (
        clk)) ;
    oai21 ix18915 (.Y (nx18914), .A0 (max_calc_comparator_first_inp2_1), .A1 (
          nx34162), .B0 (nx34165)) ;
    dff max_calc_reg_comparator_first_inp2_1 (.Q (
        max_calc_comparator_first_inp2_1), .QB (\$dummy [764]), .D (nx25433), .CLK (
        clk)) ;
    dff max_calc_reg_ans2_1 (.Q (max_calc_ans2_1), .QB (\$dummy [765]), .D (
        nx25363), .CLK (clk)) ;
    dff max_calc_reg_ans7_1 (.Q (max_calc_ans7_1), .QB (\$dummy [766]), .D (
        nx25423), .CLK (clk)) ;
    dff max_calc_reg_ans8_1 (.Q (max_calc_ans8_1), .QB (\$dummy [767]), .D (
        nx25413), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_1 (.Q (
        max_calc_comparator_first_inp1_1), .QB (nx34162), .D (nx25403), .CLK (
        clk)) ;
    dff max_calc_reg_ans1_1 (.Q (max_calc_ans1_1), .QB (\$dummy [768]), .D (
        nx25373), .CLK (clk)) ;
    dff max_calc_reg_ans6_1 (.Q (max_calc_ans6_1), .QB (\$dummy [769]), .D (
        nx25383), .CLK (clk)) ;
    dff max_calc_reg_ans5_1 (.Q (max_calc_ans5_1), .QB (\$dummy [770]), .D (
        nx25393), .CLK (clk)) ;
    oai21 ix34166 (.Y (nx34165), .A0 (nx33288), .A1 (
          max_calc_comparator_first_inp1_0), .B0 (nx18842)) ;
    xnor2 ix19141 (.Y (nx19140), .A0 (max_calc_comparator_first_inp2_15), .A1 (
          max_calc_comparator_first_inp1_15)) ;
    dff max_calc_reg_comparator_first_inp2_15 (.Q (
        max_calc_comparator_first_inp2_15), .QB (\$dummy [771]), .D (nx25553), .CLK (
        clk)) ;
    dffr labelsregfile_label2_loop1_15_fx_reg_q (.Q (label_2_output[15]), .QB (
         \$dummy [772]), .D (nx16663), .CLK (clk), .R (rst)) ;
    latch lat_label_2_input_15 (.Q (label_2_input_15), .D (nx4888), .CLK (
          nx34555)) ;
    dffr reg_label_2_input_state_machine_15 (.Q (label_2_input_state_machine_15)
         , .QB (\$dummy [773]), .D (nx15823), .CLK (clk), .R (rst)) ;
    xnor2 ix4885 (.Y (nx4884), .A0 (nx4880), .A1 (nx34182)) ;
    oai22 ix4881 (.Y (nx4880), .A0 (nx33305), .A1 (nx33477), .B0 (nx33479), .B1 (
          nx28596)) ;
    dff max_calc_reg_ans2_15 (.Q (max_calc_ans2_15), .QB (\$dummy [774]), .D (
        nx25483), .CLK (clk)) ;
    dff max_calc_reg_ans7_15 (.Q (max_calc_ans7_15), .QB (\$dummy [775]), .D (
        nx25543), .CLK (clk)) ;
    dff max_calc_reg_ans8_15 (.Q (max_calc_ans8_15), .QB (\$dummy [776]), .D (
        nx25533), .CLK (clk)) ;
    dff max_calc_reg_comparator_first_inp1_15 (.Q (
        max_calc_comparator_first_inp1_15), .QB (\$dummy [777]), .D (nx25523), .CLK (
        clk)) ;
    dffr labelsregfile_label1_loop1_15_fx_reg_q (.Q (label_1_output[15]), .QB (
         \$dummy [778]), .D (nx17513), .CLK (clk), .R (rst)) ;
    latch lat_label_1_input_15 (.Q (label_1_input_15), .D (nx6226), .CLK (
          nx34555)) ;
    dffr reg_label_1_input_state_machine_15 (.Q (label_1_input_state_machine_15)
         , .QB (\$dummy [779]), .D (nx16673), .CLK (clk), .R (rst)) ;
    xnor2 ix6223 (.Y (nx6222), .A0 (nx6218), .A1 (nx34209)) ;
    oai22 ix6219 (.Y (nx6218), .A0 (nx33503), .A1 (nx33675), .B0 (nx33677), .B1 (
          nx26636)) ;
    dff max_calc_reg_ans1_15 (.Q (max_calc_ans1_15), .QB (\$dummy [780]), .D (
        nx25493), .CLK (clk)) ;
    dff max_calc_reg_ans6_15 (.Q (max_calc_ans6_15), .QB (\$dummy [781]), .D (
        nx25503), .CLK (clk)) ;
    dff max_calc_reg_ans5_15 (.Q (max_calc_ans5_15), .QB (\$dummy [782]), .D (
        nx25513), .CLK (clk)) ;
    dffr max_calc_reg_answer_1 (.Q (answer[1]), .QB (\$dummy [783]), .D (nx25573
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_2 (.Q (answer[2]), .QB (\$dummy [784]), .D (nx25583
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_3 (.Q (answer[3]), .QB (\$dummy [785]), .D (nx25593
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_4 (.Q (answer[4]), .QB (\$dummy [786]), .D (nx25603
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_5 (.Q (answer[5]), .QB (\$dummy [787]), .D (nx25613
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_6 (.Q (answer[6]), .QB (\$dummy [788]), .D (nx25623
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_7 (.Q (answer[7]), .QB (\$dummy [789]), .D (nx25633
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_8 (.Q (answer[8]), .QB (\$dummy [790]), .D (nx25643
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_9 (.Q (answer[9]), .QB (\$dummy [791]), .D (nx25653
         ), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_10 (.Q (answer[10]), .QB (\$dummy [792]), .D (
         nx25663), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_11 (.Q (answer[11]), .QB (\$dummy [793]), .D (
         nx25673), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_12 (.Q (answer[12]), .QB (\$dummy [794]), .D (
         nx25683), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_13 (.Q (answer[13]), .QB (\$dummy [795]), .D (
         nx25693), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_14 (.Q (answer[14]), .QB (\$dummy [796]), .D (
         nx25703), .CLK (clk), .R (rst)) ;
    dffr max_calc_reg_answer_15 (.Q (answer[15]), .QB (\$dummy [797]), .D (
         nx25713), .CLK (clk), .R (rst)) ;
    tri01 tri_mdr_data_out_176 (.Y (mdr_data_out[176]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_177 (.Y (mdr_data_out[177]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_178 (.Y (mdr_data_out[178]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_179 (.Y (mdr_data_out[179]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_180 (.Y (mdr_data_out[180]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_181 (.Y (mdr_data_out[181]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_182 (.Y (mdr_data_out[182]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_183 (.Y (mdr_data_out[183]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_184 (.Y (mdr_data_out[184]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_185 (.Y (mdr_data_out[185]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_186 (.Y (mdr_data_out[186]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_187 (.Y (mdr_data_out[187]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_188 (.Y (mdr_data_out[188]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_189 (.Y (mdr_data_out[189]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_190 (.Y (mdr_data_out[190]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_191 (.Y (mdr_data_out[191]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_192 (.Y (mdr_data_out[192]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_193 (.Y (mdr_data_out[193]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_194 (.Y (mdr_data_out[194]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_195 (.Y (mdr_data_out[195]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_196 (.Y (mdr_data_out[196]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_197 (.Y (mdr_data_out[197]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_198 (.Y (mdr_data_out[198]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_199 (.Y (mdr_data_out[199]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_200 (.Y (mdr_data_out[200]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_201 (.Y (mdr_data_out[201]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_202 (.Y (mdr_data_out[202]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_203 (.Y (mdr_data_out[203]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_204 (.Y (mdr_data_out[204]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_205 (.Y (mdr_data_out[205]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_206 (.Y (mdr_data_out[206]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_207 (.Y (mdr_data_out[207]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_208 (.Y (mdr_data_out[208]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_209 (.Y (mdr_data_out[209]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_210 (.Y (mdr_data_out[210]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_211 (.Y (mdr_data_out[211]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_212 (.Y (mdr_data_out[212]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_213 (.Y (mdr_data_out[213]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_214 (.Y (mdr_data_out[214]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_215 (.Y (mdr_data_out[215]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_216 (.Y (mdr_data_out[216]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_217 (.Y (mdr_data_out[217]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_218 (.Y (mdr_data_out[218]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_219 (.Y (mdr_data_out[219]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_220 (.Y (mdr_data_out[220]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_221 (.Y (mdr_data_out[221]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_222 (.Y (mdr_data_out[222]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_223 (.Y (mdr_data_out[223]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_224 (.Y (mdr_data_out[224]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_225 (.Y (mdr_data_out[225]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_226 (.Y (mdr_data_out[226]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_227 (.Y (mdr_data_out[227]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_228 (.Y (mdr_data_out[228]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_229 (.Y (mdr_data_out[229]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_230 (.Y (mdr_data_out[230]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_231 (.Y (mdr_data_out[231]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_232 (.Y (mdr_data_out[232]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_233 (.Y (mdr_data_out[233]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_234 (.Y (mdr_data_out[234]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_235 (.Y (mdr_data_out[235]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_236 (.Y (mdr_data_out[236]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_237 (.Y (mdr_data_out[237]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_238 (.Y (mdr_data_out[238]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_239 (.Y (mdr_data_out[239]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_240 (.Y (mdr_data_out[240]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_241 (.Y (mdr_data_out[241]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_242 (.Y (mdr_data_out[242]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_243 (.Y (mdr_data_out[243]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_244 (.Y (mdr_data_out[244]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_245 (.Y (mdr_data_out[245]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_246 (.Y (mdr_data_out[246]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_247 (.Y (mdr_data_out[247]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_248 (.Y (mdr_data_out[248]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_249 (.Y (mdr_data_out[249]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_250 (.Y (mdr_data_out[250]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_251 (.Y (mdr_data_out[251]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_252 (.Y (mdr_data_out[252]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_253 (.Y (mdr_data_out[253]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_254 (.Y (mdr_data_out[254]), .A (nx25757), .E (
          initiate)) ;
    tri01 tri_mdr_data_out_255 (.Y (mdr_data_out[255]), .A (nx25757), .E (
          initiate)) ;
    dffr reg_enable_mdr_out (.Q (enable_mdr_out), .QB (\$dummy [798]), .D (
         nx25753), .CLK (clk), .R (rst)) ;
    mux21_ni ix25754 (.Y (nx25753), .A0 (enable_mdr_out), .A1 (nx190), .S0 (
             nx19296)) ;
    nor03_2x ix19297 (.Y (nx19296), .A0 (nx12895), .A1 (nx56), .A2 (nx34359)) ;
    oai21 ix34360 (.Y (nx34359), .A0 (nx25879), .A1 (nx35101), .B0 (nx868)) ;
    dffr reg_enable_mdr_in (.Q (enable_mdr_in), .QB (\$dummy [799]), .D (nx25743
         ), .CLK (clk), .R (rst)) ;
    mux21_ni ix25744 (.Y (nx25743), .A0 (nx19276), .A1 (enable_mdr_in), .S0 (
             nx34365)) ;
    nand03 ix34366 (.Y (nx34365), .A0 (nx19266), .A1 (nx26129), .A2 (nx19236)) ;
    oai21 ix19267 (.Y (nx19266), .A0 (nx34399), .A1 (nx34368), .B0 (nx174)) ;
    nor02ii ix34369 (.Y (nx34368), .A0 (nx34403), .A1 (sub_state[1])) ;
    dffr reg_enable_mar_in (.Q (enable_mar_in), .QB (\$dummy [800]), .D (nx25733
         ), .CLK (clk), .R (rst)) ;
    mux21_ni ix25734 (.Y (nx25733), .A0 (nx19250), .A1 (enable_mar_in), .S0 (
             nx34377)) ;
    ao22 ix19251 (.Y (nx19250), .A0 (nx34403), .A1 (nx174), .B0 (nx12879), .B1 (
         nx26664)) ;
    oai21 ix34378 (.Y (nx34377), .A0 (nx35157), .A1 (nx25916), .B0 (nx19240)) ;
    nor03_2x ix19233 (.Y (nx19232), .A0 (nx258), .A1 (nx12891), .A2 (nx35155)) ;
    inv01 ix19237 (.Y (nx19236), .A (nx34380)) ;
    inv01 ix15325 (.Y (nx13370), .A (nx32050)) ;
    inv01 ix15261 (.Y (nx13368), .A (nx32035)) ;
    inv01 ix15197 (.Y (nx13365), .A (nx32020)) ;
    inv01 ix15133 (.Y (nx13361), .A (nx32005)) ;
    inv01 ix15069 (.Y (nx13359), .A (nx31990)) ;
    inv01 ix15005 (.Y (nx13357), .A (nx31975)) ;
    inv01 ix14941 (.Y (nx13355), .A (nx31961)) ;
    inv01 ix31818 (.Y (nx31817), .A (nx14484)) ;
    inv01 ix31811 (.Y (nx31810), .A (nx13351)) ;
    inv01 ix14471 (.Y (nx14470), .A (nx31826)) ;
    inv01 ix31816 (.Y (nx31815), .A (nx14460)) ;
    inv01 ix14457 (.Y (nx14456), .A (nx31797)) ;
    inv01 ix31783 (.Y (nx31782), .A (nx14436)) ;
    inv01 ix31776 (.Y (nx31775), .A (nx13348)) ;
    inv01 ix14423 (.Y (nx14422), .A (nx31829)) ;
    inv01 ix31781 (.Y (nx31780), .A (nx14412)) ;
    inv01 ix14409 (.Y (nx14408), .A (nx31762)) ;
    inv01 ix31748 (.Y (nx31747), .A (nx14388)) ;
    inv01 ix31741 (.Y (nx31740), .A (nx13346)) ;
    inv01 ix14375 (.Y (nx14374), .A (nx31832)) ;
    inv01 ix31746 (.Y (nx31745), .A (nx14364)) ;
    inv01 ix14361 (.Y (nx14360), .A (nx31727)) ;
    inv01 ix31713 (.Y (nx31712), .A (nx14340)) ;
    inv01 ix31706 (.Y (nx31705), .A (nx13344)) ;
    inv01 ix14327 (.Y (nx14326), .A (nx31835)) ;
    inv01 ix31711 (.Y (nx31710), .A (nx14316)) ;
    inv01 ix14313 (.Y (nx14312), .A (nx31692)) ;
    inv01 ix31678 (.Y (nx31677), .A (nx14292)) ;
    inv01 ix31671 (.Y (nx31670), .A (nx13341)) ;
    inv01 ix14279 (.Y (nx14278), .A (nx31838)) ;
    inv01 ix31676 (.Y (nx31675), .A (nx14268)) ;
    inv01 ix14265 (.Y (nx14264), .A (nx31657)) ;
    inv01 ix31643 (.Y (nx31642), .A (nx14244)) ;
    inv01 ix31636 (.Y (nx31635), .A (nx13337)) ;
    inv01 ix14231 (.Y (nx14230), .A (nx31841)) ;
    inv01 ix31641 (.Y (nx31640), .A (nx14220)) ;
    inv01 ix14217 (.Y (nx14216), .A (nx31618)) ;
    inv01 ix31604 (.Y (nx31603), .A (nx14196)) ;
    inv01 ix31599 (.Y (nx31598), .A (nx13335)) ;
    inv01 ix14183 (.Y (nx14182), .A (nx31844)) ;
    inv01 ix14009 (.Y (nx13332), .A (nx32239)) ;
    inv01 ix13945 (.Y (nx13329), .A (nx32224)) ;
    inv01 ix13881 (.Y (nx13325), .A (nx32209)) ;
    inv01 ix13817 (.Y (nx13323), .A (nx32194)) ;
    inv01 ix13753 (.Y (nx13321), .A (nx32179)) ;
    inv01 ix13689 (.Y (nx13319), .A (nx32164)) ;
    inv01 ix13625 (.Y (nx13315), .A (nx32150)) ;
    inv01 ix31379 (.Y (nx31378), .A (nx13168)) ;
    inv01 ix31372 (.Y (nx31371), .A (nx13312)) ;
    inv01 ix13155 (.Y (nx13154), .A (nx31387)) ;
    inv01 ix31377 (.Y (nx31376), .A (nx13144)) ;
    inv01 ix13141 (.Y (nx13140), .A (nx31358)) ;
    inv01 ix31344 (.Y (nx31343), .A (nx13120)) ;
    inv01 ix31337 (.Y (nx31336), .A (nx13310)) ;
    inv01 ix13107 (.Y (nx13106), .A (nx31390)) ;
    inv01 ix31342 (.Y (nx31341), .A (nx13096)) ;
    inv01 ix13093 (.Y (nx13092), .A (nx31323)) ;
    inv01 ix31309 (.Y (nx31308), .A (nx13072)) ;
    inv01 ix31302 (.Y (nx31301), .A (nx13308)) ;
    inv01 ix13059 (.Y (nx13058), .A (nx31393)) ;
    inv01 ix31307 (.Y (nx31306), .A (nx13048)) ;
    inv01 ix13045 (.Y (nx13044), .A (nx31288)) ;
    inv01 ix31274 (.Y (nx31273), .A (nx13024)) ;
    inv01 ix31267 (.Y (nx31266), .A (nx13305)) ;
    inv01 ix13011 (.Y (nx13010), .A (nx31396)) ;
    inv01 ix31272 (.Y (nx31271), .A (nx13000)) ;
    inv01 ix12997 (.Y (nx12996), .A (nx31253)) ;
    inv01 ix31239 (.Y (nx31238), .A (nx12976)) ;
    inv01 ix31232 (.Y (nx31231), .A (nx13301)) ;
    inv01 ix12963 (.Y (nx12962), .A (nx31399)) ;
    inv01 ix31237 (.Y (nx31236), .A (nx12952)) ;
    inv01 ix12949 (.Y (nx12948), .A (nx31218)) ;
    inv01 ix31204 (.Y (nx31203), .A (nx12928)) ;
    inv01 ix31197 (.Y (nx31196), .A (nx13299)) ;
    inv01 ix12915 (.Y (nx12914), .A (nx31402)) ;
    inv01 ix31202 (.Y (nx31201), .A (nx12904)) ;
    inv01 ix12901 (.Y (nx12900), .A (nx31179)) ;
    inv01 ix31165 (.Y (nx31164), .A (nx12880)) ;
    inv01 ix31160 (.Y (nx31159), .A (nx13297)) ;
    inv01 ix12867 (.Y (nx12866), .A (nx31405)) ;
    inv01 ix12141 (.Y (nx13293), .A (nx30123)) ;
    inv01 ix12077 (.Y (nx13289), .A (nx30108)) ;
    inv01 ix12013 (.Y (nx13287), .A (nx30093)) ;
    inv01 ix11949 (.Y (nx13285), .A (nx30078)) ;
    inv01 ix11885 (.Y (nx13283), .A (nx30063)) ;
    inv01 ix11821 (.Y (nx13279), .A (nx30048)) ;
    inv01 ix11757 (.Y (nx13276), .A (nx30034)) ;
    inv01 ix29891 (.Y (nx29890), .A (nx11300)) ;
    inv01 ix29884 (.Y (nx29883), .A (nx13274)) ;
    inv01 ix11287 (.Y (nx11286), .A (nx29899)) ;
    inv01 ix29889 (.Y (nx29888), .A (nx11276)) ;
    inv01 ix11273 (.Y (nx11272), .A (nx29870)) ;
    inv01 ix29856 (.Y (nx29855), .A (nx11252)) ;
    inv01 ix29849 (.Y (nx29848), .A (nx13272)) ;
    inv01 ix11239 (.Y (nx11238), .A (nx29902)) ;
    inv01 ix29854 (.Y (nx29853), .A (nx11228)) ;
    inv01 ix11225 (.Y (nx11224), .A (nx29835)) ;
    inv01 ix29821 (.Y (nx29820), .A (nx11204)) ;
    inv01 ix29814 (.Y (nx29813), .A (nx13269)) ;
    inv01 ix11191 (.Y (nx11190), .A (nx29905)) ;
    inv01 ix29819 (.Y (nx29818), .A (nx11180)) ;
    inv01 ix11177 (.Y (nx11176), .A (nx29800)) ;
    inv01 ix29786 (.Y (nx29785), .A (nx11156)) ;
    inv01 ix29779 (.Y (nx29778), .A (nx13265)) ;
    inv01 ix11143 (.Y (nx11142), .A (nx29908)) ;
    inv01 ix29784 (.Y (nx29783), .A (nx11132)) ;
    inv01 ix11129 (.Y (nx11128), .A (nx29765)) ;
    inv01 ix29751 (.Y (nx29750), .A (nx11108)) ;
    inv01 ix29744 (.Y (nx29743), .A (nx13263)) ;
    inv01 ix11095 (.Y (nx11094), .A (nx29911)) ;
    inv01 ix29749 (.Y (nx29748), .A (nx11084)) ;
    inv01 ix11081 (.Y (nx11080), .A (nx29730)) ;
    inv01 ix29716 (.Y (nx29715), .A (nx11060)) ;
    inv01 ix29709 (.Y (nx29708), .A (nx13261)) ;
    inv01 ix11047 (.Y (nx11046), .A (nx29914)) ;
    inv01 ix29714 (.Y (nx29713), .A (nx11036)) ;
    inv01 ix11033 (.Y (nx11032), .A (nx29691)) ;
    inv01 ix29677 (.Y (nx29676), .A (nx11012)) ;
    inv01 ix29672 (.Y (nx29671), .A (nx13259)) ;
    inv01 ix10999 (.Y (nx10998), .A (nx29917)) ;
    inv01 ix10819 (.Y (nx13253), .A (nx30312)) ;
    inv01 ix10755 (.Y (nx13251), .A (nx30297)) ;
    inv01 ix10691 (.Y (nx13249), .A (nx30282)) ;
    inv01 ix10627 (.Y (nx13247), .A (nx30267)) ;
    inv01 ix10563 (.Y (nx13243), .A (nx30252)) ;
    inv01 ix10499 (.Y (nx13240), .A (nx30237)) ;
    inv01 ix10435 (.Y (nx13238), .A (nx30223)) ;
    inv01 ix29450 (.Y (nx29449), .A (nx9978)) ;
    inv01 ix29443 (.Y (nx29442), .A (nx13236)) ;
    inv01 ix9965 (.Y (nx9964), .A (nx29458)) ;
    inv01 ix29448 (.Y (nx29447), .A (nx9954)) ;
    inv01 ix9951 (.Y (nx9950), .A (nx29429)) ;
    inv01 ix29415 (.Y (nx29414), .A (nx9930)) ;
    inv01 ix29408 (.Y (nx29407), .A (nx13233)) ;
    inv01 ix9917 (.Y (nx9916), .A (nx29461)) ;
    inv01 ix29413 (.Y (nx29412), .A (nx9906)) ;
    inv01 ix9903 (.Y (nx9902), .A (nx29394)) ;
    inv01 ix29380 (.Y (nx29379), .A (nx9882)) ;
    inv01 ix29373 (.Y (nx29372), .A (nx13229)) ;
    inv01 ix9869 (.Y (nx9868), .A (nx29464)) ;
    inv01 ix29378 (.Y (nx29377), .A (nx9858)) ;
    inv01 ix9855 (.Y (nx9854), .A (nx29359)) ;
    inv01 ix29345 (.Y (nx29344), .A (nx9834)) ;
    inv01 ix29338 (.Y (nx29337), .A (nx13227)) ;
    inv01 ix9821 (.Y (nx9820), .A (nx29467)) ;
    inv01 ix29343 (.Y (nx29342), .A (nx9810)) ;
    inv01 ix9807 (.Y (nx9806), .A (nx29324)) ;
    inv01 ix29310 (.Y (nx29309), .A (nx9786)) ;
    inv01 ix29303 (.Y (nx29302), .A (nx13225)) ;
    inv01 ix9773 (.Y (nx9772), .A (nx29470)) ;
    inv01 ix29308 (.Y (nx29307), .A (nx9762)) ;
    inv01 ix9759 (.Y (nx9758), .A (nx29289)) ;
    inv01 ix29275 (.Y (nx29274), .A (nx9738)) ;
    inv01 ix29268 (.Y (nx29267), .A (nx13223)) ;
    inv01 ix9725 (.Y (nx9724), .A (nx29473)) ;
    inv01 ix29273 (.Y (nx29272), .A (nx9714)) ;
    inv01 ix9711 (.Y (nx9710), .A (nx29250)) ;
    inv01 ix29236 (.Y (nx29235), .A (nx9690)) ;
    inv01 ix29231 (.Y (nx29230), .A (nx13219)) ;
    inv01 ix9677 (.Y (nx9676), .A (nx29476)) ;
    inv01 ix9011 (.Y (nx13215), .A (nx27943)) ;
    inv01 ix8947 (.Y (nx13213), .A (nx27928)) ;
    inv01 ix8883 (.Y (nx13211), .A (nx27913)) ;
    inv01 ix8819 (.Y (nx13207), .A (nx27898)) ;
    inv01 ix8755 (.Y (nx13204), .A (nx27883)) ;
    inv01 ix8691 (.Y (nx13202), .A (nx27868)) ;
    inv01 ix8627 (.Y (nx13200), .A (nx27854)) ;
    inv01 ix8561 (.Y (nx13199), .A (nx27754)) ;
    inv01 ix8497 (.Y (nx13195), .A (nx27739)) ;
    inv01 ix8433 (.Y (nx13191), .A (nx27724)) ;
    inv01 ix8369 (.Y (nx13187), .A (nx27709)) ;
    inv01 ix8305 (.Y (nx13183), .A (nx27694)) ;
    inv01 ix8241 (.Y (nx13179), .A (nx27679)) ;
    inv01 ix8177 (.Y (nx13175), .A (nx27665)) ;
    inv01 ix27522 (.Y (nx27521), .A (nx7720)) ;
    inv01 ix27515 (.Y (nx27514), .A (nx13171)) ;
    inv01 ix7707 (.Y (nx7706), .A (nx27530)) ;
    inv01 ix27520 (.Y (nx27519), .A (nx7696)) ;
    inv01 ix7693 (.Y (nx7692), .A (nx27501)) ;
    inv01 ix27487 (.Y (nx27486), .A (nx7672)) ;
    inv01 ix27480 (.Y (nx27479), .A (nx13169)) ;
    inv01 ix7659 (.Y (nx7658), .A (nx27533)) ;
    inv01 ix27485 (.Y (nx27484), .A (nx7648)) ;
    inv01 ix7645 (.Y (nx7644), .A (nx27466)) ;
    inv01 ix27452 (.Y (nx27451), .A (nx7624)) ;
    inv01 ix27445 (.Y (nx27444), .A (nx13165)) ;
    inv01 ix7611 (.Y (nx7610), .A (nx27536)) ;
    inv01 ix27450 (.Y (nx27449), .A (nx7600)) ;
    inv01 ix7597 (.Y (nx7596), .A (nx27431)) ;
    inv01 ix27417 (.Y (nx27416), .A (nx7576)) ;
    inv01 ix27410 (.Y (nx27409), .A (nx13162)) ;
    inv01 ix7563 (.Y (nx7562), .A (nx27539)) ;
    inv01 ix27415 (.Y (nx27414), .A (nx7552)) ;
    inv01 ix7549 (.Y (nx7548), .A (nx27396)) ;
    inv01 ix27382 (.Y (nx27381), .A (nx7528)) ;
    inv01 ix27375 (.Y (nx27374), .A (nx13159)) ;
    inv01 ix7515 (.Y (nx7514), .A (nx27542)) ;
    inv01 ix27380 (.Y (nx27379), .A (nx7504)) ;
    inv01 ix7501 (.Y (nx7500), .A (nx27361)) ;
    inv01 ix27347 (.Y (nx27346), .A (nx7480)) ;
    inv01 ix27340 (.Y (nx27339), .A (nx13155)) ;
    inv01 ix7467 (.Y (nx7466), .A (nx27545)) ;
    inv01 ix27345 (.Y (nx27344), .A (nx7456)) ;
    inv01 ix7453 (.Y (nx7452), .A (nx27322)) ;
    inv01 ix27308 (.Y (nx27307), .A (nx7432)) ;
    inv01 ix27303 (.Y (nx27302), .A (nx13151)) ;
    inv01 ix7419 (.Y (nx7418), .A (nx27548)) ;
    inv01 ix27083 (.Y (nx27082), .A (nx6840)) ;
    inv01 ix27076 (.Y (nx27075), .A (nx13146)) ;
    inv01 ix6827 (.Y (nx6826), .A (nx27091)) ;
    inv01 ix27081 (.Y (nx27080), .A (nx6816)) ;
    inv01 ix6813 (.Y (nx6812), .A (nx27062)) ;
    inv01 ix27048 (.Y (nx27047), .A (nx6792)) ;
    inv01 ix27041 (.Y (nx27040), .A (nx13143)) ;
    inv01 ix6779 (.Y (nx6778), .A (nx27094)) ;
    inv01 ix27046 (.Y (nx27045), .A (nx6768)) ;
    inv01 ix6765 (.Y (nx6764), .A (nx27027)) ;
    inv01 ix27013 (.Y (nx27012), .A (nx6744)) ;
    inv01 ix27006 (.Y (nx27005), .A (nx13139)) ;
    inv01 ix6731 (.Y (nx6730), .A (nx27097)) ;
    inv01 ix27011 (.Y (nx27010), .A (nx6720)) ;
    inv01 ix6717 (.Y (nx6716), .A (nx26992)) ;
    inv01 ix26978 (.Y (nx26977), .A (nx6696)) ;
    inv01 ix26971 (.Y (nx26970), .A (nx13137)) ;
    inv01 ix6683 (.Y (nx6682), .A (nx27100)) ;
    inv01 ix26976 (.Y (nx26975), .A (nx6672)) ;
    inv01 ix6669 (.Y (nx6668), .A (nx26957)) ;
    inv01 ix26943 (.Y (nx26942), .A (nx6648)) ;
    inv01 ix26936 (.Y (nx26935), .A (nx13133)) ;
    inv01 ix6635 (.Y (nx6634), .A (nx27103)) ;
    inv01 ix26941 (.Y (nx26940), .A (nx6624)) ;
    inv01 ix6621 (.Y (nx6620), .A (nx26922)) ;
    inv01 ix26908 (.Y (nx26907), .A (nx6600)) ;
    inv01 ix26901 (.Y (nx26900), .A (nx13129)) ;
    inv01 ix6587 (.Y (nx6586), .A (nx27106)) ;
    inv01 ix26906 (.Y (nx26905), .A (nx6576)) ;
    inv01 ix6573 (.Y (nx6572), .A (nx26883)) ;
    inv01 ix26869 (.Y (nx26868), .A (nx6552)) ;
    inv01 ix26864 (.Y (nx26863), .A (nx13125)) ;
    inv01 ix6539 (.Y (nx6538), .A (nx27109)) ;
    inv01 ix6353 (.Y (nx6352), .A (nx28172)) ;
    inv01 ix6245 (.Y (nx6244), .A (nx26182)) ;
    inv01 ix6181 (.Y (nx13114), .A (nx33671)) ;
    inv01 ix6117 (.Y (nx13111), .A (nx33656)) ;
    inv01 ix6053 (.Y (nx13107), .A (nx33641)) ;
    inv01 ix5989 (.Y (nx13103), .A (nx33626)) ;
    inv01 ix5925 (.Y (nx13099), .A (nx33611)) ;
    inv01 ix5861 (.Y (nx13097), .A (nx33596)) ;
    inv01 ix5797 (.Y (nx13093), .A (nx33582)) ;
    inv01 ix26604 (.Y (nx26603), .A (nx5340)) ;
    inv01 ix26597 (.Y (nx26596), .A (nx13090)) ;
    inv01 ix5327 (.Y (nx5326), .A (nx26612)) ;
    inv01 ix26602 (.Y (nx26601), .A (nx5316)) ;
    inv01 ix5313 (.Y (nx5312), .A (nx26583)) ;
    inv01 ix26569 (.Y (nx26568), .A (nx5292)) ;
    inv01 ix26562 (.Y (nx26561), .A (nx13087)) ;
    inv01 ix5279 (.Y (nx5278), .A (nx26615)) ;
    inv01 ix26567 (.Y (nx26566), .A (nx5268)) ;
    inv01 ix5265 (.Y (nx5264), .A (nx26548)) ;
    inv01 ix26534 (.Y (nx26533), .A (nx5244)) ;
    inv01 ix26527 (.Y (nx26526), .A (nx13083)) ;
    inv01 ix5231 (.Y (nx5230), .A (nx26618)) ;
    inv01 ix26532 (.Y (nx26531), .A (nx5220)) ;
    inv01 ix5217 (.Y (nx5216), .A (nx26513)) ;
    inv01 ix26499 (.Y (nx26498), .A (nx5196)) ;
    inv01 ix26492 (.Y (nx26491), .A (nx13079)) ;
    inv01 ix5183 (.Y (nx5182), .A (nx26621)) ;
    inv01 ix26497 (.Y (nx26496), .A (nx5172)) ;
    inv01 ix5169 (.Y (nx5168), .A (nx26478)) ;
    inv01 ix26464 (.Y (nx26463), .A (nx5148)) ;
    inv01 ix26457 (.Y (nx26456), .A (nx13075)) ;
    inv01 ix5135 (.Y (nx5134), .A (nx26624)) ;
    inv01 ix26462 (.Y (nx26461), .A (nx5124)) ;
    inv01 ix5121 (.Y (nx5120), .A (nx26443)) ;
    inv01 ix26429 (.Y (nx26428), .A (nx5100)) ;
    inv01 ix26422 (.Y (nx26421), .A (nx13073)) ;
    inv01 ix5087 (.Y (nx5086), .A (nx26627)) ;
    inv01 ix26427 (.Y (nx26426), .A (nx5076)) ;
    inv01 ix5073 (.Y (nx5072), .A (nx26404)) ;
    inv01 ix26390 (.Y (nx26389), .A (nx5052)) ;
    inv01 ix26385 (.Y (nx26384), .A (nx13069)) ;
    inv01 ix5039 (.Y (nx5038), .A (nx26630)) ;
    inv01 ix4843 (.Y (nx13063), .A (nx33473)) ;
    inv01 ix4779 (.Y (nx13059), .A (nx33458)) ;
    inv01 ix4715 (.Y (nx13055), .A (nx33443)) ;
    inv01 ix4651 (.Y (nx13051), .A (nx33428)) ;
    inv01 ix4587 (.Y (nx13049), .A (nx33413)) ;
    inv01 ix4523 (.Y (nx13045), .A (nx33398)) ;
    inv01 ix4459 (.Y (nx13042), .A (nx33384)) ;
    inv01 ix28564 (.Y (nx28563), .A (nx4002)) ;
    inv01 ix28557 (.Y (nx28556), .A (nx13039)) ;
    inv01 ix3989 (.Y (nx3988), .A (nx28572)) ;
    inv01 ix28562 (.Y (nx28561), .A (nx3978)) ;
    inv01 ix3975 (.Y (nx3974), .A (nx28543)) ;
    inv01 ix28529 (.Y (nx28528), .A (nx3954)) ;
    inv01 ix28522 (.Y (nx28521), .A (nx13035)) ;
    inv01 ix3941 (.Y (nx3940), .A (nx28575)) ;
    inv01 ix28527 (.Y (nx28526), .A (nx3930)) ;
    inv01 ix3927 (.Y (nx3926), .A (nx28508)) ;
    inv01 ix28494 (.Y (nx28493), .A (nx3906)) ;
    inv01 ix28487 (.Y (nx28486), .A (nx13031)) ;
    inv01 ix3893 (.Y (nx3892), .A (nx28578)) ;
    inv01 ix28492 (.Y (nx28491), .A (nx3882)) ;
    inv01 ix3879 (.Y (nx3878), .A (nx28473)) ;
    inv01 ix28459 (.Y (nx28458), .A (nx3858)) ;
    inv01 ix28452 (.Y (nx28451), .A (nx13027)) ;
    inv01 ix3845 (.Y (nx3844), .A (nx28581)) ;
    inv01 ix28457 (.Y (nx28456), .A (nx3834)) ;
    inv01 ix3831 (.Y (nx3830), .A (nx28438)) ;
    inv01 ix28424 (.Y (nx28423), .A (nx3810)) ;
    inv01 ix28417 (.Y (nx28416), .A (nx13025)) ;
    inv01 ix3797 (.Y (nx3796), .A (nx28584)) ;
    inv01 ix28422 (.Y (nx28421), .A (nx3786)) ;
    inv01 ix3783 (.Y (nx3782), .A (nx28403)) ;
    inv01 ix28389 (.Y (nx28388), .A (nx3762)) ;
    inv01 ix28382 (.Y (nx28381), .A (nx13021)) ;
    inv01 ix3749 (.Y (nx3748), .A (nx28587)) ;
    inv01 ix28387 (.Y (nx28386), .A (nx3738)) ;
    inv01 ix3735 (.Y (nx3734), .A (nx28364)) ;
    inv01 ix28350 (.Y (nx28349), .A (nx3714)) ;
    inv01 ix28345 (.Y (nx28344), .A (nx13018)) ;
    inv01 ix3701 (.Y (nx3700), .A (nx28590)) ;
    inv01 ix3505 (.Y (nx13011), .A (nx32850)) ;
    inv01 ix3441 (.Y (nx13007), .A (nx32835)) ;
    inv01 ix3377 (.Y (nx13003), .A (nx32820)) ;
    inv01 ix3313 (.Y (nx13001), .A (nx32805)) ;
    inv01 ix3249 (.Y (nx12997), .A (nx32790)) ;
    inv01 ix3185 (.Y (nx12994), .A (nx32775)) ;
    inv01 ix3121 (.Y (nx12991), .A (nx32761)) ;
    inv01 ix29007 (.Y (nx29006), .A (nx2664)) ;
    inv01 ix29000 (.Y (nx28999), .A (nx12987)) ;
    inv01 ix2651 (.Y (nx2650), .A (nx29015)) ;
    inv01 ix29005 (.Y (nx29004), .A (nx2640)) ;
    inv01 ix2637 (.Y (nx2636), .A (nx28986)) ;
    inv01 ix28972 (.Y (nx28971), .A (nx2616)) ;
    inv01 ix28965 (.Y (nx28964), .A (nx12983)) ;
    inv01 ix2603 (.Y (nx2602), .A (nx29018)) ;
    inv01 ix28970 (.Y (nx28969), .A (nx2592)) ;
    inv01 ix2589 (.Y (nx2588), .A (nx28951)) ;
    inv01 ix28937 (.Y (nx28936), .A (nx2568)) ;
    inv01 ix28930 (.Y (nx28929), .A (nx12979)) ;
    inv01 ix2555 (.Y (nx2554), .A (nx29021)) ;
    inv01 ix28935 (.Y (nx28934), .A (nx2544)) ;
    inv01 ix2541 (.Y (nx2540), .A (nx28916)) ;
    inv01 ix28902 (.Y (nx28901), .A (nx2520)) ;
    inv01 ix28895 (.Y (nx28894), .A (nx12977)) ;
    inv01 ix2507 (.Y (nx2506), .A (nx29024)) ;
    inv01 ix28900 (.Y (nx28899), .A (nx2496)) ;
    inv01 ix2493 (.Y (nx2492), .A (nx28881)) ;
    inv01 ix28867 (.Y (nx28866), .A (nx2472)) ;
    inv01 ix28860 (.Y (nx28859), .A (nx12973)) ;
    inv01 ix2459 (.Y (nx2458), .A (nx29027)) ;
    inv01 ix28865 (.Y (nx28864), .A (nx2448)) ;
    inv01 ix2445 (.Y (nx2444), .A (nx28846)) ;
    inv01 ix28832 (.Y (nx28831), .A (nx2424)) ;
    inv01 ix28825 (.Y (nx28824), .A (nx12970)) ;
    inv01 ix2411 (.Y (nx2410), .A (nx29030)) ;
    inv01 ix28830 (.Y (nx28829), .A (nx2400)) ;
    inv01 ix2397 (.Y (nx2396), .A (nx28807)) ;
    inv01 ix28793 (.Y (nx28792), .A (nx2376)) ;
    inv01 ix28788 (.Y (nx28787), .A (nx12967)) ;
    inv01 ix2363 (.Y (nx2362), .A (nx29033)) ;
    inv01 ix2167 (.Y (nx12959), .A (nx32654)) ;
    inv01 ix2103 (.Y (nx12955), .A (nx32639)) ;
    inv01 ix2039 (.Y (nx12953), .A (nx32624)) ;
    inv01 ix1975 (.Y (nx12949), .A (nx32609)) ;
    inv01 ix1911 (.Y (nx12946), .A (nx32594)) ;
    inv01 ix1847 (.Y (nx12943), .A (nx32579)) ;
    inv01 ix1783 (.Y (nx12939), .A (nx32565)) ;
    inv01 ix30936 (.Y (nx30935), .A (nx1326)) ;
    inv01 ix30929 (.Y (nx30928), .A (nx12935)) ;
    inv01 ix1313 (.Y (nx1312), .A (nx30944)) ;
    inv01 ix30934 (.Y (nx30933), .A (nx1302)) ;
    inv01 ix1299 (.Y (nx1298), .A (nx30915)) ;
    inv01 ix30901 (.Y (nx30900), .A (nx1278)) ;
    inv01 ix30894 (.Y (nx30893), .A (nx12931)) ;
    inv01 ix1265 (.Y (nx1264), .A (nx30947)) ;
    inv01 ix30899 (.Y (nx30898), .A (nx1254)) ;
    inv01 ix1251 (.Y (nx1250), .A (nx30880)) ;
    inv01 ix30866 (.Y (nx30865), .A (nx1230)) ;
    inv01 ix30859 (.Y (nx30858), .A (nx12929)) ;
    inv01 ix1217 (.Y (nx1216), .A (nx30950)) ;
    inv01 ix30864 (.Y (nx30863), .A (nx1206)) ;
    inv01 ix1203 (.Y (nx1202), .A (nx30845)) ;
    inv01 ix30831 (.Y (nx30830), .A (nx1182)) ;
    inv01 ix30824 (.Y (nx30823), .A (nx12925)) ;
    inv01 ix1169 (.Y (nx1168), .A (nx30953)) ;
    inv01 ix30829 (.Y (nx30828), .A (nx1158)) ;
    inv01 ix1155 (.Y (nx1154), .A (nx30810)) ;
    inv01 ix30796 (.Y (nx30795), .A (nx1134)) ;
    inv01 ix30789 (.Y (nx30788), .A (nx12922)) ;
    inv01 ix1121 (.Y (nx1120), .A (nx30956)) ;
    inv01 ix30794 (.Y (nx30793), .A (nx1110)) ;
    inv01 ix1107 (.Y (nx1106), .A (nx30775)) ;
    inv01 ix30761 (.Y (nx30760), .A (nx1086)) ;
    inv01 ix30754 (.Y (nx30753), .A (nx12919)) ;
    inv01 ix1073 (.Y (nx1072), .A (nx30959)) ;
    inv01 ix30759 (.Y (nx30758), .A (nx1062)) ;
    inv01 ix1059 (.Y (nx1058), .A (nx30736)) ;
    inv01 ix30722 (.Y (nx30721), .A (nx1038)) ;
    inv01 ix30717 (.Y (nx30716), .A (nx12915)) ;
    inv01 ix1025 (.Y (nx1024), .A (nx30962)) ;
    inv01 ix657 (.Y (nx656), .A (nx26056)) ;
    inv01 ix549 (.Y (nx548), .A (nx26001)) ;
    inv01 ix25836 (.Y (nx25835), .A (nx516)) ;
    inv01 ix457 (.Y (nx12898), .A (nx25962)) ;
    inv01 ix25920 (.Y (nx25919), .A (nx334)) ;
    inv01 ix853 (.Y (nx12895), .A (nx26129)) ;
    inv01 ix187 (.Y (nx186), .A (nx25907)) ;
    inv01 ix25917 (.Y (nx25916), .A (nx174)) ;
    inv01 ix25814 (.Y (nx25813), .A (nx12891)) ;
    inv01 ix26665 (.Y (nx26664), .A (nx38)) ;
    inv01 ix49 (.Y (nx12885), .A (nx25944)) ;
    inv01 ix25901 (.Y (nx25900), .A (nx12879)) ;
    inv02 ix34388 (.Y (nx34389), .A (nx35783)) ;
    inv02 ix34390 (.Y (nx34391), .A (nx35783)) ;
    inv02 ix34392 (.Y (nx34393), .A (nx35779)) ;
    inv02 ix34394 (.Y (nx34395), .A (nx35779)) ;
    inv02 ix34396 (.Y (nx34397), .A (nx35791)) ;
    inv02 ix34398 (.Y (nx34399), .A (nx35791)) ;
    buf02 ix34400 (.Y (nx34401), .A (sub_state[0])) ;
    buf02 ix34402 (.Y (nx34403), .A (sub_state[0])) ;
    inv02 ix34404 (.Y (nx34405), .A (nx35153)) ;
    inv02 ix34406 (.Y (nx34407), .A (nx35153)) ;
    inv02 ix34408 (.Y (nx34409), .A (nx35919)) ;
    inv02 ix34418 (.Y (nx34419), .A (nx35925)) ;
    inv02 ix34428 (.Y (nx34429), .A (nx35925)) ;
    inv02 ix34456 (.Y (nx34457), .A (ready_signal)) ;
    inv02 ix34458 (.Y (nx34459), .A (nx35589)) ;
    inv02 ix34460 (.Y (nx34461), .A (nx35589)) ;
    inv02 ix34462 (.Y (nx34463), .A (nx35589)) ;
    inv02 ix34464 (.Y (nx34465), .A (nx35589)) ;
    inv02 ix34466 (.Y (nx34467), .A (nx35589)) ;
    inv02 ix34468 (.Y (nx34469), .A (nx35591)) ;
    inv02 ix34470 (.Y (nx34471), .A (nx35591)) ;
    inv02 ix34472 (.Y (nx34473), .A (nx35591)) ;
    inv02 ix34474 (.Y (nx34475), .A (nx35591)) ;
    inv02 ix34476 (.Y (nx34477), .A (nx35591)) ;
    inv02 ix34478 (.Y (nx34479), .A (nx35591)) ;
    inv02 ix34480 (.Y (nx34481), .A (nx35591)) ;
    inv02 ix34482 (.Y (nx34483), .A (nx35593)) ;
    inv02 ix34484 (.Y (nx34485), .A (nx35593)) ;
    inv02 ix34486 (.Y (nx34487), .A (nx35593)) ;
    inv02 ix34488 (.Y (nx34489), .A (nx35593)) ;
    inv02 ix34490 (.Y (nx34491), .A (nx35593)) ;
    inv02 ix34492 (.Y (nx34493), .A (nx35593)) ;
    inv02 ix34494 (.Y (nx34495), .A (nx35101)) ;
    inv02 ix34498 (.Y (nx34499), .A (nx25999)) ;
    inv02 ix34500 (.Y (nx34501), .A (nx35799)) ;
    buf02 ix34502 (.Y (nx34503), .A (enable_address)) ;
    buf02 ix34504 (.Y (nx34505), .A (enable_address)) ;
    buf02 ix34506 (.Y (nx34507), .A (nx350)) ;
    buf02 ix34508 (.Y (nx34509), .A (nx350)) ;
    inv02 ix34510 (.Y (nx34511), .A (nx35263)) ;
    inv02 ix34512 (.Y (nx34513), .A (nx35265)) ;
    inv02 ix34514 (.Y (nx34515), .A (nx35265)) ;
    inv02 ix34516 (.Y (nx34517), .A (nx35265)) ;
    inv02 ix34518 (.Y (nx34519), .A (nx35265)) ;
    inv02 ix34520 (.Y (nx34521), .A (nx35265)) ;
    inv02 ix34522 (.Y (nx34523), .A (nx35265)) ;
    inv02 ix34524 (.Y (nx34525), .A (nx35265)) ;
    inv02 ix34526 (.Y (nx34527), .A (nx35267)) ;
    inv02 ix34528 (.Y (nx34529), .A (nx35267)) ;
    inv02 ix34530 (.Y (nx34531), .A (nx35267)) ;
    inv02 ix34532 (.Y (nx34533), .A (nx35267)) ;
    inv02 ix34534 (.Y (nx34535), .A (nx35267)) ;
    inv02 ix34536 (.Y (nx34537), .A (nx35267)) ;
    inv02 ix34538 (.Y (nx34539), .A (nx35267)) ;
    inv02 ix34540 (.Y (nx34541), .A (nx35269)) ;
    inv02 ix34542 (.Y (nx34543), .A (nx35269)) ;
    inv02 ix34544 (.Y (nx34545), .A (nx35269)) ;
    inv02 ix34546 (.Y (nx34547), .A (nx35269)) ;
    inv02 ix34548 (.Y (nx34549), .A (nx35269)) ;
    inv02 ix34550 (.Y (nx34551), .A (nx35269)) ;
    inv02 ix34552 (.Y (nx34553), .A (nx35269)) ;
    inv02 ix34554 (.Y (nx34555), .A (nx35271)) ;
    inv02 ix34556 (.Y (nx34557), .A (nx36147)) ;
    inv02 ix34570 (.Y (nx34571), .A (nx36155)) ;
    inv02 ix34578 (.Y (nx34579), .A (nx30744)) ;
    inv02 ix34580 (.Y (nx34581), .A (nx30744)) ;
    inv02 ix34582 (.Y (nx34583), .A (nx30744)) ;
    inv02 ix34588 (.Y (nx34589), .A (nx36093)) ;
    inv02 ix34602 (.Y (nx34603), .A (nx36101)) ;
    inv02 ix34610 (.Y (nx34611), .A (nx28815)) ;
    inv02 ix34612 (.Y (nx34613), .A (nx28815)) ;
    inv02 ix34614 (.Y (nx34615), .A (nx28815)) ;
    inv02 ix34620 (.Y (nx34621), .A (nx36077)) ;
    inv02 ix34634 (.Y (nx34635), .A (nx36085)) ;
    inv02 ix34642 (.Y (nx34643), .A (nx28372)) ;
    inv02 ix34644 (.Y (nx34645), .A (nx28372)) ;
    inv02 ix34646 (.Y (nx34647), .A (nx28372)) ;
    inv02 ix34652 (.Y (nx34653), .A (nx36003)) ;
    inv02 ix34666 (.Y (nx34667), .A (nx36011)) ;
    inv02 ix34674 (.Y (nx34675), .A (nx26412)) ;
    inv02 ix34676 (.Y (nx34677), .A (nx26412)) ;
    inv02 ix34678 (.Y (nx34679), .A (nx26412)) ;
    inv02 ix34704 (.Y (nx34705), .A (nx35977)) ;
    inv02 ix34736 (.Y (nx34737), .A (nx34735)) ;
    inv02 ix34738 (.Y (nx34739), .A (nx35843)) ;
    inv02 ix34740 (.Y (nx34741), .A (nx35843)) ;
    inv02 ix34742 (.Y (nx34743), .A (nx35843)) ;
    inv02 ix34744 (.Y (nx34745), .A (nx35843)) ;
    inv02 ix34746 (.Y (nx34747), .A (nx35361)) ;
    inv02 ix34748 (.Y (nx34749), .A (nx35361)) ;
    inv02 ix34750 (.Y (nx34751), .A (nx35361)) ;
    inv02 ix34752 (.Y (nx34753), .A (nx36063)) ;
    inv02 ix34754 (.Y (nx34755), .A (nx36063)) ;
    inv02 ix34756 (.Y (nx34757), .A (nx36063)) ;
    inv02 ix34758 (.Y (nx34759), .A (nx36063)) ;
    inv02 ix34760 (.Y (nx34761), .A (nx36063)) ;
    inv02 ix34762 (.Y (nx34763), .A (nx36063)) ;
    inv02 ix34764 (.Y (nx34765), .A (nx36063)) ;
    inv02 ix34766 (.Y (nx34767), .A (nx36067)) ;
    inv02 ix34768 (.Y (nx34769), .A (nx36067)) ;
    inv02 ix34770 (.Y (nx34771), .A (nx36067)) ;
    inv02 ix34772 (.Y (nx34773), .A (nx36067)) ;
    inv02 ix34774 (.Y (nx34775), .A (nx36067)) ;
    inv02 ix34776 (.Y (nx34777), .A (nx36067)) ;
    inv02 ix34778 (.Y (nx34779), .A (nx36067)) ;
    inv02 ix34780 (.Y (nx34781), .A (nx36071)) ;
    inv02 ix34782 (.Y (nx34783), .A (nx36071)) ;
    inv02 ix34784 (.Y (nx34785), .A (nx36071)) ;
    inv02 ix34786 (.Y (nx34787), .A (nx36071)) ;
    inv02 ix34788 (.Y (nx34789), .A (nx36071)) ;
    inv02 ix34790 (.Y (nx34791), .A (nx36071)) ;
    inv02 ix34792 (.Y (nx34793), .A (nx36071)) ;
    inv02 ix34794 (.Y (nx34795), .A (nx36075)) ;
    inv02 ix34796 (.Y (nx34797), .A (nx36075)) ;
    inv02 ix34798 (.Y (nx34799), .A (nx36075)) ;
    inv02 ix34800 (.Y (nx34801), .A (nx36075)) ;
    inv02 ix34802 (.Y (nx34803), .A (nx36075)) ;
    inv02 ix34804 (.Y (nx34805), .A (nx36075)) ;
    inv02 ix34806 (.Y (nx34807), .A (nx36075)) ;
    inv02 ix34808 (.Y (nx34809), .A (nx35371)) ;
    inv02 ix34810 (.Y (nx34811), .A (nx35371)) ;
    inv02 ix34812 (.Y (nx34813), .A (nx35371)) ;
    inv02 ix34814 (.Y (nx34815), .A (nx35371)) ;
    inv02 ix34816 (.Y (nx34817), .A (nx35371)) ;
    inv02 ix34818 (.Y (nx34819), .A (nx35371)) ;
    inv02 ix34832 (.Y (nx34833), .A (nx36031)) ;
    inv02 ix34846 (.Y (nx34847), .A (nx36039)) ;
    inv02 ix34854 (.Y (nx34855), .A (nx26891)) ;
    inv02 ix34856 (.Y (nx34857), .A (nx26891)) ;
    inv02 ix34858 (.Y (nx34859), .A (nx26891)) ;
    inv02 ix34864 (.Y (nx34865), .A (nx36047)) ;
    inv02 ix34878 (.Y (nx34879), .A (nx36055)) ;
    inv02 ix34886 (.Y (nx34887), .A (nx27330)) ;
    inv02 ix34888 (.Y (nx34889), .A (nx27330)) ;
    inv02 ix34890 (.Y (nx34891), .A (nx27330)) ;
    inv02 ix34924 (.Y (nx34925), .A (nx36109)) ;
    inv02 ix34938 (.Y (nx34939), .A (nx36117)) ;
    inv02 ix34946 (.Y (nx34947), .A (nx29258)) ;
    inv02 ix34948 (.Y (nx34949), .A (nx29258)) ;
    inv02 ix34950 (.Y (nx34951), .A (nx29258)) ;
    inv02 ix34956 (.Y (nx34957), .A (nx36131)) ;
    inv02 ix34970 (.Y (nx34971), .A (nx36139)) ;
    inv02 ix34978 (.Y (nx34979), .A (nx29699)) ;
    inv02 ix34980 (.Y (nx34981), .A (nx29699)) ;
    inv02 ix34982 (.Y (nx34983), .A (nx29699)) ;
    inv02 ix34996 (.Y (nx34997), .A (nx36163)) ;
    inv02 ix35010 (.Y (nx35011), .A (nx36171)) ;
    inv02 ix35018 (.Y (nx35019), .A (nx31187)) ;
    inv02 ix35020 (.Y (nx35021), .A (nx31187)) ;
    inv02 ix35022 (.Y (nx35023), .A (nx31187)) ;
    inv02 ix35028 (.Y (nx35029), .A (nx36179)) ;
    inv02 ix35042 (.Y (nx35043), .A (nx36187)) ;
    inv02 ix35050 (.Y (nx35051), .A (nx31626)) ;
    inv02 ix35052 (.Y (nx35053), .A (nx31626)) ;
    inv02 ix35054 (.Y (nx35055), .A (nx31626)) ;
    buf02 ix35094 (.Y (nx35095), .A (nx25827)) ;
    buf02 ix35096 (.Y (nx35097), .A (nx25827)) ;
    inv02 ix35098 (.Y (nx35099), .A (nx12893)) ;
    inv02 ix35100 (.Y (nx35101), .A (nx12893)) ;
    inv02 ix35102 (.Y (nx35103), .A (nx36201)) ;
    inv02 ix35148 (.Y (nx35149), .A (nx4)) ;
    inv02 ix35152 (.Y (nx35153), .A (nx35713)) ;
    inv02 ix35154 (.Y (nx35155), .A (nx12882)) ;
    buf02 ix35156 (.Y (nx35157), .A (nx25896)) ;
    buf02 ix35158 (.Y (nx35159), .A (nx25937)) ;
    buf02 ix35160 (.Y (nx35161), .A (nx25937)) ;
    inv02 ix35162 (.Y (nx35163), .A (enable_decoder_dst_booth)) ;
    inv02 ix35164 (.Y (nx35165), .A (nx36307)) ;
    inv02 ix35166 (.Y (nx35167), .A (nx36307)) ;
    inv02 ix35168 (.Y (nx35169), .A (nx36307)) ;
    inv02 ix35170 (.Y (nx35171), .A (nx36307)) ;
    inv02 ix35172 (.Y (nx35173), .A (max_calc_state_2)) ;
    inv02 ix35174 (.Y (nx35175), .A (nx36299)) ;
    inv02 ix35176 (.Y (nx35177), .A (nx36299)) ;
    inv02 ix35178 (.Y (nx35179), .A (nx36299)) ;
    inv02 ix35180 (.Y (nx35181), .A (nx36299)) ;
    inv02 ix35182 (.Y (nx35183), .A (nx36299)) ;
    inv02 ix35184 (.Y (nx35185), .A (nx36299)) ;
    inv02 ix35186 (.Y (nx35187), .A (max_calc_state_1)) ;
    inv02 ix35188 (.Y (nx35189), .A (nx36331)) ;
    inv02 ix35190 (.Y (nx35191), .A (nx36331)) ;
    inv02 ix35192 (.Y (nx35193), .A (
          booth_booth_integrtaion_0_shift_reg_output_9)) ;
    inv02 ix35194 (.Y (nx35195), .A (nx36327)) ;
    inv02 ix35196 (.Y (nx35197), .A (nx36327)) ;
    inv02 ix35198 (.Y (nx35199), .A (nx36327)) ;
    inv01 ix35200 (.Y (nx35201), .A (
          booth_booth_integrtaion_0_shift_reg_output_0)) ;
    buf02 ix35204 (.Y (nx35205), .A (nx26386)) ;
    buf02 ix35206 (.Y (nx35207), .A (nx26423)) ;
    buf02 ix35208 (.Y (nx35209), .A (nx26458)) ;
    buf02 ix35210 (.Y (nx35211), .A (nx26493)) ;
    buf02 ix35212 (.Y (nx35213), .A (nx26528)) ;
    buf02 ix35214 (.Y (nx35215), .A (nx26563)) ;
    buf02 ix35216 (.Y (nx35217), .A (nx26598)) ;
    inv02 ix35262 (.Y (nx35263), .A (nx36277)) ;
    inv02 ix35264 (.Y (nx35265), .A (nx36277)) ;
    inv02 ix35266 (.Y (nx35267), .A (nx36277)) ;
    inv02 ix35268 (.Y (nx35269), .A (nx36277)) ;
    inv02 ix35270 (.Y (nx35271), .A (nx36277)) ;
    inv02 ix35300 (.Y (nx35301), .A (
          booth_booth_integrtaion_8_shift_reg_output_9)) ;
    inv02 ix35302 (.Y (nx35303), .A (nx36341)) ;
    inv02 ix35304 (.Y (nx35305), .A (nx36341)) ;
    inv02 ix35306 (.Y (nx35307), .A (nx36341)) ;
    inv01 ix35308 (.Y (nx35309), .A (
          booth_booth_integrtaion_8_shift_reg_output_0)) ;
    buf02 ix35312 (.Y (nx35313), .A (nx26865)) ;
    buf02 ix35314 (.Y (nx35315), .A (nx26902)) ;
    buf02 ix35316 (.Y (nx35317), .A (nx26937)) ;
    buf02 ix35318 (.Y (nx35319), .A (nx26972)) ;
    buf02 ix35320 (.Y (nx35321), .A (nx27007)) ;
    buf02 ix35322 (.Y (nx35323), .A (nx27042)) ;
    buf02 ix35324 (.Y (nx35325), .A (nx27077)) ;
    inv02 ix35326 (.Y (nx35327), .A (
          booth_booth_integrtaion_9_shift_reg_output_9)) ;
    inv02 ix35328 (.Y (nx35329), .A (nx36345)) ;
    inv02 ix35330 (.Y (nx35331), .A (nx36345)) ;
    inv02 ix35332 (.Y (nx35333), .A (nx36345)) ;
    inv01 ix35334 (.Y (nx35335), .A (
          booth_booth_integrtaion_9_shift_reg_output_0)) ;
    buf02 ix35338 (.Y (nx35339), .A (nx27304)) ;
    buf02 ix35340 (.Y (nx35341), .A (nx27341)) ;
    buf02 ix35342 (.Y (nx35343), .A (nx27376)) ;
    buf02 ix35344 (.Y (nx35345), .A (nx27411)) ;
    buf02 ix35346 (.Y (nx35347), .A (nx27446)) ;
    buf02 ix35348 (.Y (nx35349), .A (nx27481)) ;
    buf02 ix35350 (.Y (nx35351), .A (nx27516)) ;
    inv02 ix35360 (.Y (nx35361), .A (nx36281)) ;
    inv02 ix35362 (.Y (nx35363), .A (nx36337)) ;
    inv02 ix35364 (.Y (nx35365), .A (nx36337)) ;
    inv02 ix35366 (.Y (nx35367), .A (nx36337)) ;
    inv02 ix35368 (.Y (nx35369), .A (nx36337)) ;
    inv02 ix35370 (.Y (nx35371), .A (nx36337)) ;
    inv02 ix35372 (.Y (nx35373), .A (
          booth_booth_integrtaion_1_shift_reg_output_9)) ;
    inv02 ix35374 (.Y (nx35375), .A (nx36323)) ;
    inv02 ix35376 (.Y (nx35377), .A (nx36323)) ;
    inv02 ix35378 (.Y (nx35379), .A (nx36323)) ;
    inv01 ix35380 (.Y (nx35381), .A (
          booth_booth_integrtaion_1_shift_reg_output_0)) ;
    buf02 ix35384 (.Y (nx35385), .A (nx28346)) ;
    buf02 ix35386 (.Y (nx35387), .A (nx28383)) ;
    buf02 ix35388 (.Y (nx35389), .A (nx28418)) ;
    buf02 ix35390 (.Y (nx35391), .A (nx28453)) ;
    buf02 ix35392 (.Y (nx35393), .A (nx28488)) ;
    buf02 ix35394 (.Y (nx35395), .A (nx28523)) ;
    buf02 ix35396 (.Y (nx35397), .A (nx28558)) ;
    inv02 ix35398 (.Y (nx35399), .A (
          booth_booth_integrtaion_2_shift_reg_output_9)) ;
    inv02 ix35400 (.Y (nx35401), .A (nx36319)) ;
    inv02 ix35402 (.Y (nx35403), .A (nx36319)) ;
    inv02 ix35404 (.Y (nx35405), .A (nx36319)) ;
    inv01 ix35406 (.Y (nx35407), .A (
          booth_booth_integrtaion_2_shift_reg_output_0)) ;
    buf02 ix35410 (.Y (nx35411), .A (nx28789)) ;
    buf02 ix35412 (.Y (nx35413), .A (nx28826)) ;
    buf02 ix35414 (.Y (nx35415), .A (nx28861)) ;
    buf02 ix35416 (.Y (nx35417), .A (nx28896)) ;
    buf02 ix35418 (.Y (nx35419), .A (nx28931)) ;
    buf02 ix35420 (.Y (nx35421), .A (nx28966)) ;
    buf02 ix35422 (.Y (nx35423), .A (nx29001)) ;
    inv02 ix35424 (.Y (nx35425), .A (
          booth_booth_integrtaion_4_shift_reg_output_9)) ;
    inv02 ix35426 (.Y (nx35427), .A (nx36349)) ;
    inv02 ix35428 (.Y (nx35429), .A (nx36349)) ;
    inv02 ix35430 (.Y (nx35431), .A (nx36349)) ;
    inv01 ix35432 (.Y (nx35433), .A (
          booth_booth_integrtaion_4_shift_reg_output_0)) ;
    buf02 ix35436 (.Y (nx35437), .A (nx29232)) ;
    buf02 ix35438 (.Y (nx35439), .A (nx29269)) ;
    buf02 ix35440 (.Y (nx35441), .A (nx29304)) ;
    buf02 ix35442 (.Y (nx35443), .A (nx29339)) ;
    buf02 ix35444 (.Y (nx35445), .A (nx29374)) ;
    buf02 ix35446 (.Y (nx35447), .A (nx29409)) ;
    buf02 ix35448 (.Y (nx35449), .A (nx29444)) ;
    inv02 ix35452 (.Y (nx35453), .A (nx36195)) ;
    inv02 ix35454 (.Y (nx35455), .A (nx36195)) ;
    inv02 ix35456 (.Y (nx35457), .A (nx36195)) ;
    inv02 ix35458 (.Y (nx35459), .A (nx36195)) ;
    inv02 ix35460 (.Y (nx35461), .A (nx36195)) ;
    inv02 ix35462 (.Y (nx35463), .A (nx36125)) ;
    inv02 ix35464 (.Y (nx35465), .A (nx36125)) ;
    inv02 ix35466 (.Y (nx35467), .A (nx36125)) ;
    inv02 ix35468 (.Y (nx35469), .A (nx36125)) ;
    inv02 ix35472 (.Y (nx35473), .A (
          booth_booth_integrtaion_5_shift_reg_output_9)) ;
    inv02 ix35474 (.Y (nx35475), .A (nx36353)) ;
    inv02 ix35476 (.Y (nx35477), .A (nx36353)) ;
    inv02 ix35478 (.Y (nx35479), .A (nx36353)) ;
    inv01 ix35480 (.Y (nx35481), .A (
          booth_booth_integrtaion_5_shift_reg_output_0)) ;
    buf02 ix35484 (.Y (nx35485), .A (nx29673)) ;
    buf02 ix35486 (.Y (nx35487), .A (nx29710)) ;
    buf02 ix35488 (.Y (nx35489), .A (nx29745)) ;
    buf02 ix35490 (.Y (nx35491), .A (nx29780)) ;
    buf02 ix35492 (.Y (nx35493), .A (nx29815)) ;
    buf02 ix35494 (.Y (nx35495), .A (nx29850)) ;
    buf02 ix35496 (.Y (nx35497), .A (nx29885)) ;
    inv02 ix35498 (.Y (nx35499), .A (
          booth_booth_integrtaion_3_shift_reg_output_9)) ;
    inv02 ix35500 (.Y (nx35501), .A (nx36315)) ;
    inv02 ix35502 (.Y (nx35503), .A (nx36315)) ;
    inv02 ix35504 (.Y (nx35505), .A (nx36315)) ;
    inv01 ix35506 (.Y (nx35507), .A (
          booth_booth_integrtaion_3_shift_reg_output_0)) ;
    buf02 ix35510 (.Y (nx35511), .A (nx30718)) ;
    buf02 ix35512 (.Y (nx35513), .A (nx30755)) ;
    buf02 ix35514 (.Y (nx35515), .A (nx30790)) ;
    buf02 ix35516 (.Y (nx35517), .A (nx30825)) ;
    buf02 ix35518 (.Y (nx35519), .A (nx30860)) ;
    buf02 ix35520 (.Y (nx35521), .A (nx30895)) ;
    buf02 ix35522 (.Y (nx35523), .A (nx30930)) ;
    inv02 ix35524 (.Y (nx35525), .A (
          booth_booth_integrtaion_6_shift_reg_output_9)) ;
    inv02 ix35526 (.Y (nx35527), .A (nx36357)) ;
    inv02 ix35528 (.Y (nx35529), .A (nx36357)) ;
    inv02 ix35530 (.Y (nx35531), .A (nx36357)) ;
    inv01 ix35532 (.Y (nx35533), .A (
          booth_booth_integrtaion_6_shift_reg_output_0)) ;
    buf02 ix35536 (.Y (nx35537), .A (nx31161)) ;
    buf02 ix35538 (.Y (nx35539), .A (nx31198)) ;
    buf02 ix35540 (.Y (nx35541), .A (nx31233)) ;
    buf02 ix35542 (.Y (nx35543), .A (nx31268)) ;
    buf02 ix35544 (.Y (nx35545), .A (nx31303)) ;
    buf02 ix35546 (.Y (nx35547), .A (nx31338)) ;
    buf02 ix35548 (.Y (nx35549), .A (nx31373)) ;
    inv02 ix35550 (.Y (nx35551), .A (
          booth_booth_integrtaion_7_shift_reg_output_9)) ;
    inv02 ix35552 (.Y (nx35553), .A (nx36361)) ;
    inv02 ix35554 (.Y (nx35555), .A (nx36361)) ;
    inv02 ix35556 (.Y (nx35557), .A (nx36361)) ;
    inv01 ix35558 (.Y (nx35559), .A (
          booth_booth_integrtaion_7_shift_reg_output_0)) ;
    buf02 ix35562 (.Y (nx35563), .A (nx31600)) ;
    buf02 ix35564 (.Y (nx35565), .A (nx31637)) ;
    buf02 ix35566 (.Y (nx35567), .A (nx31672)) ;
    buf02 ix35568 (.Y (nx35569), .A (nx31707)) ;
    buf02 ix35570 (.Y (nx35571), .A (nx31742)) ;
    buf02 ix35572 (.Y (nx35573), .A (nx31777)) ;
    buf02 ix35574 (.Y (nx35575), .A (nx31812)) ;
    inv02 ix35588 (.Y (nx35589), .A (nx34457)) ;
    inv02 ix35590 (.Y (nx35591), .A (nx34457)) ;
    inv02 ix35592 (.Y (nx35593), .A (nx34457)) ;
    inv02 ix35594 (.Y (nx35595), .A (nx25854)) ;
    inv02 ix35596 (.Y (nx35597), .A (nx36365)) ;
    inv02 ix35598 (.Y (nx35599), .A (nx36365)) ;
    inv02 ix35600 (.Y (nx35601), .A (nx36365)) ;
    inv02 ix35602 (.Y (nx35603), .A (nx26669)) ;
    inv02 ix35604 (.Y (nx35605), .A (nx36373)) ;
    inv02 ix35606 (.Y (nx35607), .A (nx36373)) ;
    inv02 ix35608 (.Y (nx35609), .A (nx36373)) ;
    inv02 ix35614 (.Y (nx35615), .A (ready_signal)) ;
    nand02 ix13624 (.Y (nx13623), .A0 (nx35911), .A1 (nx35919)) ;
    mux21_ni ix13614 (.Y (nx13613), .A0 (nx34409), .A1 (
             booth_shift_Reg_adder_0_output_17), .S0 (nx35911)) ;
    mux21_ni ix13604 (.Y (nx13603), .A0 (booth_shift_Reg_adder_0_output_17), .A1 (
             booth_shift_Reg_adder_0_output_16), .S0 (nx35911)) ;
    mux21_ni ix13594 (.Y (nx13593), .A0 (booth_shift_Reg_adder_0_output_16), .A1 (
             booth_shift_Reg_adder_0_output_15), .S0 (nx35911)) ;
    mux21_ni ix13584 (.Y (nx13583), .A0 (booth_shift_Reg_adder_0_output_15), .A1 (
             booth_shift_Reg_adder_0_output_14), .S0 (nx35911)) ;
    mux21_ni ix13574 (.Y (nx13573), .A0 (booth_shift_Reg_adder_0_output_14), .A1 (
             booth_shift_Reg_adder_0_output_13), .S0 (nx35911)) ;
    mux21_ni ix13564 (.Y (nx13563), .A0 (booth_shift_Reg_adder_0_output_13), .A1 (
             booth_shift_Reg_adder_0_output_12), .S0 (nx35911)) ;
    mux21_ni ix13554 (.Y (nx13553), .A0 (booth_shift_Reg_adder_0_output_12), .A1 (
             booth_shift_Reg_adder_0_output_11), .S0 (nx35913)) ;
    mux21_ni ix13544 (.Y (nx13543), .A0 (booth_shift_Reg_adder_0_output_11), .A1 (
             booth_shift_Reg_adder_0_output_10), .S0 (nx35913)) ;
    mux21_ni ix13534 (.Y (nx13533), .A0 (booth_shift_Reg_adder_0_output_10), .A1 (
             booth_shift_Reg_adder_0_output_9), .S0 (nx35913)) ;
    mux21_ni ix13524 (.Y (nx13523), .A0 (booth_shift_Reg_adder_0_output_9), .A1 (
             booth_shift_Reg_adder_0_output_8), .S0 (nx35913)) ;
    mux21_ni ix13514 (.Y (nx13513), .A0 (booth_shift_Reg_adder_0_output_8), .A1 (
             booth_shift_Reg_adder_0_output_7), .S0 (nx35913)) ;
    mux21_ni ix13504 (.Y (nx13503), .A0 (booth_shift_Reg_adder_0_output_7), .A1 (
             booth_shift_Reg_adder_0_output_6), .S0 (nx35913)) ;
    mux21_ni ix13494 (.Y (nx13493), .A0 (booth_shift_Reg_adder_0_output_6), .A1 (
             booth_shift_Reg_adder_0_output_5), .S0 (nx35913)) ;
    mux21_ni ix13484 (.Y (nx13483), .A0 (booth_shift_Reg_adder_0_output_5), .A1 (
             booth_shift_Reg_adder_0_output_4), .S0 (nx35915)) ;
    mux21_ni ix13474 (.Y (nx13473), .A0 (booth_shift_Reg_adder_0_output_4), .A1 (
             booth_shift_Reg_adder_0_output_3), .S0 (nx35915)) ;
    mux21_ni ix13464 (.Y (nx13463), .A0 (booth_shift_Reg_adder_0_output_3), .A1 (
             booth_shift_Reg_adder_0_output_2), .S0 (nx35915)) ;
    mux21_ni ix13454 (.Y (nx13453), .A0 (booth_shift_Reg_adder_0_output_2), .A1 (
             booth_shift_Reg_adder_0_output_1), .S0 (nx35915)) ;
    mux21_ni ix13444 (.Y (nx13443), .A0 (booth_shift_Reg_adder_0_output_1), .A1 (
             booth_shift_Reg_adder_0_output_0), .S0 (nx35915)) ;
    nor02ii ix13430 (.Y (nx13429), .A0 (nx35915), .A1 (
            booth_shift_Reg_adder_0_output_0)) ;
    mux21 ix13424 (.Y (nx13423), .A0 (nx34457), .A1 (nx35153), .S0 (nx64)) ;
    ao221 ix831 (.Y (nx830), .A0 (nx35791), .A1 (nx172), .B0 (nx25944), .B1 (
          nx35713), .C0 (nx35621)) ;
    ao32 ix13634 (.Y (nx13633), .A0 (nx35783), .A1 (nx35779), .A2 (nx25907), .B0 (
         sub_state[2]), .B1 (nx35623)) ;
    inv01 ix35622 (.Y (nx35623), .A (nx12883)) ;
    nand02 ix14094 (.Y (nx14093), .A0 (nx35783), .A1 (nx25832)) ;
    mux21_ni ix13834 (.Y (nx13833), .A0 (num_in_2), .A1 (num_out_2), .S0 (
             nx35795)) ;
    ao22 ix497 (.Y (nx496), .A0 (mdr_data_out[2]), .A1 (nx12893), .B0 (nx35625)
         , .B1 (nx35713)) ;
    inv01 ix35624 (.Y (nx35625), .A (nx25821)) ;
    mux21 ix13664 (.Y (nx13663), .A0 (nx35153), .A1 (nx35799), .S0 (nx35097)) ;
    mux21_ni ix13714 (.Y (nx13713), .A0 (num_in_0), .A1 (num_out_0), .S0 (
             nx35795)) ;
    ao22 ix377 (.Y (nx376), .A0 (mdr_data_out[0]), .A1 (nx12893), .B0 (nx35627)
         , .B1 (nx35713)) ;
    inv01 ix35626 (.Y (nx35627), .A (nx25864)) ;
    and03 ix805 (.Y (nx12879), .A0 (nx25857), .A1 (nx35783), .A2 (state[1])) ;
    and03 ix173 (.Y (nx172), .A0 (state[0]), .A1 (nx35783), .A2 (nx35779)) ;
    nor03_2x ix25860 (.Y (nx4), .A0 (nx25857), .A1 (state[2]), .A2 (nx35779)) ;
    ao21 ix811 (.Y (nx12877), .A0 (nx25857), .A1 (nx35779), .B0 (nx35783)) ;
    xor2 ix25865 (.Y (nx25864), .A0 (alu_inp1_0), .A1 (nx25935)) ;
    mux21_ni ix391 (.Y (nx390), .A0 (address_out_0), .A1 (num_out_0), .S0 (
             nx35713)) ;
    nor02ii ix25875 (.Y (nx25874), .A0 (sub_state[1]), .A1 (nx12893)) ;
    nor02ii ix27 (.Y (nx26), .A0 (nx25879), .A1 (nx12887)) ;
    ao32 ix21 (.Y (nx20), .A0 (nx12887), .A1 (nx35791), .A2 (nx35629), .B0 (
         nx25944), .B1 (nx35713)) ;
    inv01 ix35628 (.Y (nx35629), .A (nx34401)) ;
    and02 ix175 (.Y (nx174), .A0 (nx35785), .A1 (nx35779)) ;
    nand02 ix25890 (.Y (nx12882), .A0 (nx35915), .A1 (nx35589)) ;
    nor02ii ix25894 (.Y (nx25893), .A0 (nx174), .A1 (nx35153)) ;
    ao32 ix335 (.Y (nx334), .A0 (nx35631), .A1 (nx35791), .A2 (nx320), .B0 (
         nx35101), .B1 (nx25907)) ;
    nand02 ix25906 (.Y (nx35631), .A0 (nx186), .A1 (nx172)) ;
    nor02ii ix25908 (.Y (nx25907), .A0 (nx35157), .A1 (nx35791)) ;
    and03 ix225 (.Y (nx12893), .A0 (nx25857), .A1 (nx35785), .A2 (nx35781)) ;
    mux21 ix243 (.Y (nx242), .A0 (nx35793), .A1 (nx35153), .S0 (nx35101)) ;
    mux21_ni ix13774 (.Y (nx13773), .A0 (num_in_1), .A1 (num_out_1), .S0 (
             nx35795)) ;
    mux21_ni ix413 (.Y (nx412), .A0 (alu_inp1_0), .A1 (nx34499), .S0 (nx25935)
             ) ;
    xor2 ix25963 (.Y (nx25962), .A0 (alu_inp1_1), .A1 (nx35799)) ;
    mux21_ni ix449 (.Y (nx448), .A0 (address_out_1), .A1 (num_out_1), .S0 (
             nx35713)) ;
    mux21_ni ix13884 (.Y (nx13883), .A0 (num_in_3), .A1 (num_out_3), .S0 (
             nx35795)) ;
    xnor2 ix25987 (.Y (nx25986), .A0 (nx25998), .A1 (nx35799)) ;
    mux21_ni ix481 (.Y (nx480), .A0 (address_out_2), .A1 (num_out_2), .S0 (
             nx35715)) ;
    xor2 ix26002 (.Y (nx26001), .A0 (alu_inp1_3), .A1 (nx35801)) ;
    mux21_ni ix541 (.Y (nx540), .A0 (address_out_3), .A1 (num_out_3), .S0 (
             nx35715)) ;
    mux21_ni ix13934 (.Y (nx13933), .A0 (num_in_4), .A1 (num_out_4), .S0 (
             nx35795)) ;
    ao22 ix607 (.Y (nx606), .A0 (mdr_data_out[4]), .A1 (nx12893), .B0 (nx35633)
         , .B1 (nx35715)) ;
    inv01 ix35632 (.Y (nx35633), .A (nx26022)) ;
    xnor2 ix26028 (.Y (nx26027), .A0 (nx26039), .A1 (nx35801)) ;
    mux21_ni ix591 (.Y (nx590), .A0 (address_out_4), .A1 (num_out_4), .S0 (
             nx35715)) ;
    or04 ix26045 (.Y (nx26044), .A0 (num_out_5), .A1 (num_out_6), .A2 (num_out_7
         ), .A3 (nx35917)) ;
    mux21 ix13984 (.Y (nx13983), .A0 (nx26069), .A1 (nx26046), .S0 (nx35795)) ;
    xor2 ix26057 (.Y (nx26056), .A0 (alu_inp1_5), .A1 (nx35801)) ;
    mux21_ni ix649 (.Y (nx648), .A0 (address_out_5), .A1 (num_out_5), .S0 (
             nx35715)) ;
    mux21_ni ix14034 (.Y (nx14033), .A0 (num_in_6), .A1 (num_out_6), .S0 (
             nx35797)) ;
    ao22 ix715 (.Y (nx714), .A0 (mdr_data_out[6]), .A1 (nx12893), .B0 (nx35635)
         , .B1 (nx35715)) ;
    inv01 ix35634 (.Y (nx35635), .A (nx26078)) ;
    xnor2 ix26084 (.Y (nx26083), .A0 (nx26095), .A1 (nx35801)) ;
    mux21_ni ix699 (.Y (nx698), .A0 (address_out_6), .A1 (num_out_6), .S0 (
             nx35715)) ;
    mux21 ix14084 (.Y (nx14083), .A0 (nx26122), .A1 (nx26099), .S0 (nx35797)) ;
    xor2 ix26110 (.Y (nx26109), .A0 (alu_inp1_7), .A1 (nx35801)) ;
    mux21_ni ix755 (.Y (nx754), .A0 (address_out_7), .A1 (num_out_7), .S0 (
             nx35717)) ;
    and03 ix843 (.Y (nx12909), .A0 (nx25857), .A1 (state[2]), .A2 (nx35781)) ;
    oai21 ix26140 (.Y (nx35621), .A0 (nx35793), .A1 (nx35101), .B0 (nx35637)) ;
    or04 ix819 (.Y (nx35637), .A0 (nx12891), .A1 (nx25900), .A2 (nx35155), .A3 (
         nx35157)) ;
    and04 ix65 (.Y (nx64), .A0 (nx35785), .A1 (state[1]), .A2 (nx35639), .A3 (
          nx25942)) ;
    inv01 ix35638 (.Y (nx35639), .A (nx56)) ;
    or02 ix26183 (.Y (nx26182), .A0 (nx26176), .A1 (max_calc_start)) ;
    and02 ix26192 (.Y (nx26191), .A0 (nx26176), .A1 (nx26180)) ;
    xnor2 ix26195 (.Y (nx26194), .A0 (nx26188), .A1 (nx35977)) ;
    ao32 ix17554 (.Y (nx17553), .A0 (nx35641), .A1 (nx26203), .A2 (
         max_calc_start), .B0 (nx36331), .B1 (nx26191)) ;
    inv01 ix35640 (.Y (nx35641), .A (nx26194)) ;
    ao22 ix17564 (.Y (nx17563), .A0 (max_calc_start), .A1 (nx35843), .B0 (
         max_calc_state_3), .B1 (nx26191)) ;
    nor03_2x ix6277 (.Y (nx34735), .A0 (nx26188), .A1 (nx35977), .A2 (nx35643)
             ) ;
    inv01 ix35642 (.Y (nx35643), .A (nx26201)) ;
    and02 ix26202 (.Y (nx26201), .A0 (nx36299), .A1 (nx26203)) ;
    mux21_ni ix25564 (.Y (nx25563), .A0 (answer[0]), .A1 (nx13121), .S0 (nx35741
             )) ;
    mux21_ni ix19151 (.Y (nx13121), .A0 (max_calc_comparator_first_inp2_0), .A1 (
             max_calc_comparator_first_inp1_0), .S0 (nx35905)) ;
    mux21_ni ix19634 (.Y (nx19633), .A0 (max_calc_comparator_first_inp1_0), .A1 (
             nx9512), .S0 (nx36281)) ;
    mux21_ni ix9513 (.Y (nx9512), .A0 (nx9508), .A1 (nx6388), .S0 (nx35959)) ;
    mux21_ni ix6389 (.Y (nx6388), .A0 (max_calc_ans1_0), .A1 (label_1_output[0])
             , .S0 (nx35977)) ;
    mux21_ni ix17224 (.Y (nx17223), .A0 (label_1_output[0]), .A1 (
             label_1_input_0), .S0 (nx36241)) ;
    mux21_ni ix17214 (.Y (nx17213), .A0 (label_1_input_state_machine_0), .A1 (
             mdr_data_out[0]), .S0 (nx36201)) ;
    mux21_ni ix17204 (.Y (nx17203), .A0 (nx35731), .A1 (nx5736), .S0 (nx35199)
             ) ;
    mux21_ni ix5737 (.Y (nx5736), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_0_1), .S0 (nx36011)) ;
    mux21_ni ix17194 (.Y (nx17193), .A0 (booth_booth_integration_output_0_1), .A1 (
             nx5724), .S0 (nx35199)) ;
    mux21_ni ix5725 (.Y (nx5724), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_0_2), .S0 (nx36011)) ;
    mux21_ni ix17184 (.Y (nx17183), .A0 (booth_booth_integration_output_0_2), .A1 (
             nx5712), .S0 (nx35199)) ;
    mux21_ni ix5713 (.Y (nx5712), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_0_3), .S0 (nx36011)) ;
    mux21_ni ix17174 (.Y (nx17173), .A0 (booth_booth_integration_output_0_3), .A1 (
             nx5700), .S0 (nx35199)) ;
    mux21_ni ix5701 (.Y (nx5700), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_0_4), .S0 (nx36011)) ;
    mux21_ni ix17164 (.Y (nx17163), .A0 (booth_booth_integration_output_0_4), .A1 (
             nx5688), .S0 (nx35199)) ;
    mux21_ni ix5689 (.Y (nx5688), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_0_5), .S0 (nx36011)) ;
    mux21_ni ix17154 (.Y (nx17153), .A0 (booth_booth_integration_output_0_5), .A1 (
             nx5676), .S0 (nx35199)) ;
    mux21_ni ix5677 (.Y (nx5676), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_0_6), .S0 (nx36013)) ;
    mux21_ni ix17144 (.Y (nx17143), .A0 (booth_booth_integration_output_0_6), .A1 (
             nx5664), .S0 (nx35199)) ;
    mux21_ni ix5665 (.Y (nx5664), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_0_7), .S0 (nx36013)) ;
    mux21_ni ix17134 (.Y (nx17133), .A0 (booth_booth_integration_output_0_7), .A1 (
             nx5652), .S0 (nx36003)) ;
    mux21_ni ix5653 (.Y (nx5652), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_0_8), .S0 (nx36013)) ;
    mux21_ni ix17124 (.Y (nx17123), .A0 (booth_booth_integration_output_0_8), .A1 (
             nx5640), .S0 (nx36003)) ;
    mux21_ni ix5641 (.Y (nx5640), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_0_9), .S0 (nx36013)) ;
    mux21_ni ix17114 (.Y (nx17113), .A0 (booth_booth_integration_output_0_9), .A1 (
             nx5628), .S0 (nx36003)) ;
    mux21_ni ix5629 (.Y (nx5628), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_0_10), .S0 (nx36013)) ;
    mux21_ni ix17104 (.Y (nx17103), .A0 (booth_booth_integration_output_0_10), .A1 (
             nx5616), .S0 (nx36005)) ;
    mux21_ni ix5617 (.Y (nx5616), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_0_11), .S0 (nx36013)) ;
    mux21_ni ix17094 (.Y (nx17093), .A0 (booth_booth_integration_output_0_11), .A1 (
             nx5604), .S0 (nx36005)) ;
    mux21_ni ix5605 (.Y (nx5604), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_0_12), .S0 (nx36013)) ;
    mux21_ni ix17084 (.Y (nx17083), .A0 (booth_booth_integration_output_0_12), .A1 (
             nx5592), .S0 (nx36005)) ;
    mux21_ni ix5593 (.Y (nx5592), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_0_13), .S0 (nx36015)) ;
    mux21_ni ix17074 (.Y (nx17073), .A0 (booth_booth_integration_output_0_13), .A1 (
             nx5580), .S0 (nx36005)) ;
    mux21_ni ix5581 (.Y (nx5580), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_0_14), .S0 (nx36015)) ;
    mux21_ni ix17064 (.Y (nx17063), .A0 (booth_booth_integration_output_0_14), .A1 (
             nx5568), .S0 (nx36005)) ;
    mux21_ni ix5569 (.Y (nx5568), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_0_15), .S0 (nx36015)) ;
    mux21 ix17054 (.Y (nx17053), .A0 (nx26634), .A1 (nx26276), .S0 (nx36005)) ;
    mux21_ni ix16704 (.Y (nx16703), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_0), .A1 (nx34667), .S0 (
             nx35803)) ;
    and02 ix16690 (.Y (nx16689), .A0 (nx36327), .A1 (
          booth_booth_integrtaion_0_shift_Reg_count_0)) ;
    mux21_ni ix16884 (.Y (nx16883), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_9), .A1 (nx34653), .S0 (
             nx35803)) ;
    mux21_ni ix16874 (.Y (nx16873), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_8), .S0 (nx36005)) ;
    mux21_ni ix16864 (.Y (nx16863), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_8), .S0 (nx35803)) ;
    mux21_ni ix16854 (.Y (nx16853), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_7), .S0 (nx36007)) ;
    mux21_ni ix16844 (.Y (nx16843), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_7), .S0 (nx35803)) ;
    mux21_ni ix16834 (.Y (nx16833), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_6), .S0 (nx36007)) ;
    mux21_ni ix16824 (.Y (nx16823), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_6), .S0 (nx35803)) ;
    mux21_ni ix16814 (.Y (nx16813), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_5), .S0 (nx36007)) ;
    mux21_ni ix16804 (.Y (nx16803), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_5), .S0 (nx35803)) ;
    mux21_ni ix16794 (.Y (nx16793), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_4), .S0 (nx36007)) ;
    mux21_ni ix16784 (.Y (nx16783), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_4), .S0 (nx35805)) ;
    mux21_ni ix16774 (.Y (nx16773), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_3), .S0 (nx36007)) ;
    mux21_ni ix16764 (.Y (nx16763), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_3), .S0 (nx35805)) ;
    mux21_ni ix16754 (.Y (nx16753), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_2), .S0 (nx36007)) ;
    mux21_ni ix16744 (.Y (nx16743), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_2), .S0 (nx35805)) ;
    mux21_ni ix16734 (.Y (nx16733), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_1), .S0 (nx36007)) ;
    mux21_ni ix16724 (.Y (nx16723), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_0_shift_Reg_output_1), .S0 (nx35805)) ;
    mux21_ni ix16714 (.Y (nx16713), .A0 (
             booth_booth_integrtaion_0_shift_Reg_count_1), .A1 (nx34667), .S0 (
             nx36009)) ;
    and02 ix5009 (.Y (nx5008), .A0 (nx26349), .A1 (nx35731)) ;
    or03 ix26352 (.Y (nx26351), .A0 (nx26353), .A1 (
         booth_booth_integrtaion_0_shift_reg_output_0), .A2 (nx36327)) ;
    mux21_ni ix17044 (.Y (nx17043), .A0 (
             booth_booth_integrtaion_0_booth_output_16), .A1 (nx5538), .S0 (
             nx36009)) ;
    nor02ii ix5539 (.Y (nx5538), .A0 (nx26360), .A1 (nx36015)) ;
    nor02ii ix5015 (.Y (nx5014), .A0 (nx26344), .A1 (
            booth_booth_integrtaion_0_booth_output_16)) ;
    xor2 ix5533 (.Y (nx13067), .A0 (nx26366), .A1 (nx26630)) ;
    xor2 ix5521 (.Y (nx13069), .A0 (nx26391), .A1 (nx35205)) ;
    mux21_ni ix17024 (.Y (nx17023), .A0 (
             booth_booth_integrtaion_0_booth_output_18), .A1 (nx5514), .S0 (
             nx36009)) ;
    nor02ii ix5515 (.Y (nx5514), .A0 (nx26381), .A1 (nx36015)) ;
    xor2 ix5509 (.Y (nx13071), .A0 (nx26396), .A1 (nx26627)) ;
    or02 ix26413 (.Y (nx26412), .A0 (nx26349), .A1 (nx35733)) ;
    xor2 ix5497 (.Y (nx13073), .A0 (nx26430), .A1 (nx35207)) ;
    mux21_ni ix17004 (.Y (nx17003), .A0 (
             booth_booth_integrtaion_0_booth_output_20), .A1 (nx5490), .S0 (
             nx36009)) ;
    nor02ii ix5491 (.Y (nx5490), .A0 (nx26418), .A1 (nx36015)) ;
    xor2 ix5485 (.Y (nx13074), .A0 (nx26435), .A1 (nx26624)) ;
    xor2 ix5473 (.Y (nx13075), .A0 (nx26465), .A1 (nx35209)) ;
    mux21_ni ix16984 (.Y (nx16983), .A0 (
             booth_booth_integrtaion_0_booth_output_22), .A1 (nx5466), .S0 (
             nx36009)) ;
    nor02ii ix5467 (.Y (nx5466), .A0 (nx26453), .A1 (nx36015)) ;
    xor2 ix5461 (.Y (nx13077), .A0 (nx26470), .A1 (nx26621)) ;
    xor2 ix5449 (.Y (nx13079), .A0 (nx26500), .A1 (nx35211)) ;
    mux21_ni ix16964 (.Y (nx16963), .A0 (
             booth_booth_integrtaion_0_booth_output_24), .A1 (nx5442), .S0 (
             nx36009)) ;
    nor02ii ix5443 (.Y (nx5442), .A0 (nx26488), .A1 (nx36017)) ;
    xor2 ix5437 (.Y (nx13081), .A0 (nx26505), .A1 (nx26618)) ;
    xor2 ix5425 (.Y (nx13083), .A0 (nx26535), .A1 (nx35213)) ;
    mux21_ni ix16944 (.Y (nx16943), .A0 (
             booth_booth_integrtaion_0_booth_output_26), .A1 (nx5418), .S0 (
             nx36009)) ;
    nor02ii ix5419 (.Y (nx5418), .A0 (nx26523), .A1 (nx36017)) ;
    xor2 ix5413 (.Y (nx13085), .A0 (nx26540), .A1 (nx26615)) ;
    xor2 ix5401 (.Y (nx13087), .A0 (nx26570), .A1 (nx35215)) ;
    mux21_ni ix16924 (.Y (nx16923), .A0 (
             booth_booth_integrtaion_0_booth_output_28), .A1 (nx5394), .S0 (
             nx35197)) ;
    nor02ii ix5395 (.Y (nx5394), .A0 (nx26558), .A1 (nx36017)) ;
    xor2 ix5389 (.Y (nx13089), .A0 (nx26575), .A1 (nx26612)) ;
    xor2 ix5377 (.Y (nx13090), .A0 (nx26605), .A1 (nx35217)) ;
    mux21_ni ix16904 (.Y (nx16903), .A0 (
             booth_booth_integrtaion_0_booth_output_31), .A1 (nx5370), .S0 (
             nx35197)) ;
    nor02ii ix5371 (.Y (nx5370), .A0 (nx26593), .A1 (nx36017)) ;
    xor2 ix5365 (.Y (nx5364), .A0 (nx26605), .A1 (nx26608)) ;
    nor02ii ix5551 (.Y (nx5550), .A0 (nx5014), .A1 (nx36017)) ;
    oai21 ix26658 (.Y (nx846), .A0 (nx35781), .A1 (nx25857), .B0 (nx35785)) ;
    and02 ix26667 (.Y (nx26666), .A0 (nx35791), .A1 (sub_state[1])) ;
    nor02ii ix26670 (.Y (nx26669), .A0 (sel_dst_0), .A1 (nx35919)) ;
    mux21_ni ix17584 (.Y (nx17583), .A0 (nx13121), .A1 (max_calc_ans1_0), .S0 (
             nx35851)) ;
    nand03 ix6379 (.Y (nx34821), .A0 (nx35959), .A1 (nx26203), .A2 (nx36291)) ;
    mux21_ni ix9509 (.Y (nx9508), .A0 (max_calc_ans5_0), .A1 (max_calc_ans6_0), 
             .S0 (nx35977)) ;
    mux21_ni ix17594 (.Y (nx17593), .A0 (max_calc_ans6_0), .A1 (nx13121), .S0 (
             nx36021)) ;
    nor02ii ix26683 (.Y (nx35289), .A0 (nx36381), .A1 (nx26194)) ;
    mux21_ni ix19624 (.Y (nx19623), .A0 (max_calc_ans5_0), .A1 (nx9498), .S0 (
             nx36291)) ;
    mux21 ix9499 (.Y (nx9498), .A0 (nx27133), .A1 (nx26693), .S0 (nx35861)) ;
    mux21_ni ix18144 (.Y (nx18143), .A0 (label_9_output[0]), .A1 (
             label_9_input_0), .S0 (nx36241)) ;
    mux21_ni ix18134 (.Y (nx18133), .A0 (label_9_input_state_machine_0), .A1 (
             mdr_data_out[128]), .S0 (nx36201)) ;
    mux21_ni ix18124 (.Y (nx18123), .A0 (nx35755), .A1 (nx7236), .S0 (nx35307)
             ) ;
    mux21_ni ix7237 (.Y (nx7236), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_8_1), .S0 (nx36039)) ;
    mux21_ni ix18114 (.Y (nx18113), .A0 (booth_booth_integration_output_8_1), .A1 (
             nx7224), .S0 (nx35307)) ;
    mux21_ni ix7225 (.Y (nx7224), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_8_2), .S0 (nx36039)) ;
    mux21_ni ix18104 (.Y (nx18103), .A0 (booth_booth_integration_output_8_2), .A1 (
             nx7212), .S0 (nx35307)) ;
    mux21_ni ix7213 (.Y (nx7212), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_8_3), .S0 (nx36039)) ;
    mux21_ni ix18094 (.Y (nx18093), .A0 (booth_booth_integration_output_8_3), .A1 (
             nx7200), .S0 (nx35307)) ;
    mux21_ni ix7201 (.Y (nx7200), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_8_4), .S0 (nx36039)) ;
    mux21_ni ix18084 (.Y (nx18083), .A0 (booth_booth_integration_output_8_4), .A1 (
             nx7188), .S0 (nx35307)) ;
    mux21_ni ix7189 (.Y (nx7188), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_8_5), .S0 (nx36039)) ;
    mux21_ni ix18074 (.Y (nx18073), .A0 (booth_booth_integration_output_8_5), .A1 (
             nx7176), .S0 (nx35307)) ;
    mux21_ni ix7177 (.Y (nx7176), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_8_6), .S0 (nx36041)) ;
    mux21_ni ix18064 (.Y (nx18063), .A0 (booth_booth_integration_output_8_6), .A1 (
             nx7164), .S0 (nx35307)) ;
    mux21_ni ix7165 (.Y (nx7164), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_8_7), .S0 (nx36041)) ;
    mux21_ni ix18054 (.Y (nx18053), .A0 (booth_booth_integration_output_8_7), .A1 (
             nx7152), .S0 (nx36031)) ;
    mux21_ni ix7153 (.Y (nx7152), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_8_8), .S0 (nx36041)) ;
    mux21_ni ix18044 (.Y (nx18043), .A0 (booth_booth_integration_output_8_8), .A1 (
             nx7140), .S0 (nx36031)) ;
    mux21_ni ix7141 (.Y (nx7140), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_8_9), .S0 (nx36041)) ;
    mux21_ni ix18034 (.Y (nx18033), .A0 (booth_booth_integration_output_8_9), .A1 (
             nx7128), .S0 (nx36031)) ;
    mux21_ni ix7129 (.Y (nx7128), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_8_10), .S0 (nx36041)) ;
    mux21_ni ix18024 (.Y (nx18023), .A0 (booth_booth_integration_output_8_10), .A1 (
             nx7116), .S0 (nx36033)) ;
    mux21_ni ix7117 (.Y (nx7116), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_8_11), .S0 (nx36041)) ;
    mux21_ni ix18014 (.Y (nx18013), .A0 (booth_booth_integration_output_8_11), .A1 (
             nx7104), .S0 (nx36033)) ;
    mux21_ni ix7105 (.Y (nx7104), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_8_12), .S0 (nx36041)) ;
    mux21_ni ix18004 (.Y (nx18003), .A0 (booth_booth_integration_output_8_12), .A1 (
             nx7092), .S0 (nx36033)) ;
    mux21_ni ix7093 (.Y (nx7092), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_8_13), .S0 (nx36043)) ;
    mux21_ni ix17994 (.Y (nx17993), .A0 (booth_booth_integration_output_8_13), .A1 (
             nx7080), .S0 (nx36033)) ;
    mux21_ni ix7081 (.Y (nx7080), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_8_14), .S0 (nx36043)) ;
    mux21_ni ix17984 (.Y (nx17983), .A0 (booth_booth_integration_output_8_14), .A1 (
             nx7068), .S0 (nx36033)) ;
    mux21_ni ix7069 (.Y (nx7068), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_8_15), .S0 (nx36043)) ;
    mux21 ix17974 (.Y (nx17973), .A0 (nx27113), .A1 (nx26755), .S0 (nx36033)) ;
    mux21_ni ix17624 (.Y (nx17623), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_0), .A1 (nx34847), .S0 (
             nx35807)) ;
    and02 ix17610 (.Y (nx17609), .A0 (nx36341), .A1 (
          booth_booth_integrtaion_8_shift_Reg_count_0)) ;
    mux21_ni ix17804 (.Y (nx17803), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_9), .A1 (nx34833), .S0 (
             nx35807)) ;
    mux21_ni ix17794 (.Y (nx17793), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_8), .S0 (nx36033)) ;
    mux21_ni ix17784 (.Y (nx17783), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_8), .S0 (nx35807)) ;
    mux21_ni ix17774 (.Y (nx17773), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_7), .S0 (nx36035)) ;
    mux21_ni ix17764 (.Y (nx17763), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_7), .S0 (nx35807)) ;
    mux21_ni ix17754 (.Y (nx17753), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_6), .S0 (nx36035)) ;
    mux21_ni ix17744 (.Y (nx17743), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_6), .S0 (nx35807)) ;
    mux21_ni ix17734 (.Y (nx17733), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_5), .S0 (nx36035)) ;
    mux21_ni ix17724 (.Y (nx17723), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_5), .S0 (nx35807)) ;
    mux21_ni ix17714 (.Y (nx17713), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_4), .S0 (nx36035)) ;
    mux21_ni ix17704 (.Y (nx17703), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_4), .S0 (nx35809)) ;
    mux21_ni ix17694 (.Y (nx17693), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_3), .S0 (nx36035)) ;
    mux21_ni ix17684 (.Y (nx17683), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_3), .S0 (nx35809)) ;
    mux21_ni ix17674 (.Y (nx17673), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_2), .S0 (nx36035)) ;
    mux21_ni ix17664 (.Y (nx17663), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_2), .S0 (nx35809)) ;
    mux21_ni ix17654 (.Y (nx17653), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_1), .S0 (nx36035)) ;
    mux21_ni ix17644 (.Y (nx17643), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_8_shift_Reg_output_1), .S0 (nx35809)) ;
    mux21_ni ix17634 (.Y (nx17633), .A0 (
             booth_booth_integrtaion_8_shift_Reg_count_1), .A1 (nx34847), .S0 (
             nx36037)) ;
    and02 ix6509 (.Y (nx6508), .A0 (nx26828), .A1 (nx35755)) ;
    or03 ix26831 (.Y (nx26830), .A0 (nx26832), .A1 (
         booth_booth_integrtaion_8_shift_reg_output_0), .A2 (nx36341)) ;
    mux21_ni ix17964 (.Y (nx17963), .A0 (
             booth_booth_integrtaion_8_booth_output_16), .A1 (nx7038), .S0 (
             nx36037)) ;
    nor02ii ix7039 (.Y (nx7038), .A0 (nx26839), .A1 (nx36043)) ;
    nor02ii ix6515 (.Y (nx6514), .A0 (nx26823), .A1 (
            booth_booth_integrtaion_8_booth_output_16)) ;
    xor2 ix7033 (.Y (nx13123), .A0 (nx26845), .A1 (nx27109)) ;
    xor2 ix7021 (.Y (nx13125), .A0 (nx26870), .A1 (nx35313)) ;
    mux21_ni ix17944 (.Y (nx17943), .A0 (
             booth_booth_integrtaion_8_booth_output_18), .A1 (nx7014), .S0 (
             nx36037)) ;
    nor02ii ix7015 (.Y (nx7014), .A0 (nx26860), .A1 (nx36043)) ;
    xor2 ix7009 (.Y (nx13127), .A0 (nx26875), .A1 (nx27106)) ;
    or02 ix26892 (.Y (nx26891), .A0 (nx26828), .A1 (nx35757)) ;
    xor2 ix6997 (.Y (nx13129), .A0 (nx26909), .A1 (nx35315)) ;
    mux21_ni ix17924 (.Y (nx17923), .A0 (
             booth_booth_integrtaion_8_booth_output_20), .A1 (nx6990), .S0 (
             nx36037)) ;
    nor02ii ix6991 (.Y (nx6990), .A0 (nx26897), .A1 (nx36043)) ;
    xor2 ix6985 (.Y (nx13131), .A0 (nx26914), .A1 (nx27103)) ;
    xor2 ix6973 (.Y (nx13133), .A0 (nx26944), .A1 (nx35317)) ;
    mux21_ni ix17904 (.Y (nx17903), .A0 (
             booth_booth_integrtaion_8_booth_output_22), .A1 (nx6966), .S0 (
             nx36037)) ;
    nor02ii ix6967 (.Y (nx6966), .A0 (nx26932), .A1 (nx36043)) ;
    xor2 ix6961 (.Y (nx13135), .A0 (nx26949), .A1 (nx27100)) ;
    xor2 ix6949 (.Y (nx13137), .A0 (nx26979), .A1 (nx35319)) ;
    mux21_ni ix17884 (.Y (nx17883), .A0 (
             booth_booth_integrtaion_8_booth_output_24), .A1 (nx6942), .S0 (
             nx36037)) ;
    nor02ii ix6943 (.Y (nx6942), .A0 (nx26967), .A1 (nx36045)) ;
    xor2 ix6937 (.Y (nx13138), .A0 (nx26984), .A1 (nx27097)) ;
    xor2 ix6925 (.Y (nx13139), .A0 (nx27014), .A1 (nx35321)) ;
    mux21_ni ix17864 (.Y (nx17863), .A0 (
             booth_booth_integrtaion_8_booth_output_26), .A1 (nx6918), .S0 (
             nx36037)) ;
    nor02ii ix6919 (.Y (nx6918), .A0 (nx27002), .A1 (nx36045)) ;
    xor2 ix6913 (.Y (nx13141), .A0 (nx27019), .A1 (nx27094)) ;
    xor2 ix6901 (.Y (nx13143), .A0 (nx27049), .A1 (nx35323)) ;
    mux21_ni ix17844 (.Y (nx17843), .A0 (
             booth_booth_integrtaion_8_booth_output_28), .A1 (nx6894), .S0 (
             nx35305)) ;
    nor02ii ix6895 (.Y (nx6894), .A0 (nx27037), .A1 (nx36045)) ;
    xor2 ix6889 (.Y (nx13145), .A0 (nx27054), .A1 (nx27091)) ;
    xor2 ix6877 (.Y (nx13146), .A0 (nx27084), .A1 (nx35325)) ;
    mux21_ni ix17824 (.Y (nx17823), .A0 (
             booth_booth_integrtaion_8_booth_output_31), .A1 (nx6870), .S0 (
             nx35305)) ;
    nor02ii ix6871 (.Y (nx6870), .A0 (nx27072), .A1 (nx36045)) ;
    xor2 ix6865 (.Y (nx6864), .A0 (nx27084), .A1 (nx27087)) ;
    nor02ii ix7051 (.Y (nx7050), .A0 (nx6514), .A1 (nx36045)) ;
    mux21_ni ix18714 (.Y (nx18713), .A0 (label_10_output[0]), .A1 (
             label_10_input_0), .S0 (nx36241)) ;
    mux21_ni ix18704 (.Y (nx18703), .A0 (label_10_input_state_machine_0), .A1 (
             mdr_data_out[144]), .S0 (nx36201)) ;
    mux21_ni ix18694 (.Y (nx18693), .A0 (nx35759), .A1 (nx8116), .S0 (nx35333)
             ) ;
    mux21_ni ix8117 (.Y (nx8116), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_9_1), .S0 (nx36055)) ;
    mux21_ni ix18684 (.Y (nx18683), .A0 (booth_booth_integration_output_9_1), .A1 (
             nx8104), .S0 (nx35333)) ;
    mux21_ni ix8105 (.Y (nx8104), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_9_2), .S0 (nx36055)) ;
    mux21_ni ix18674 (.Y (nx18673), .A0 (booth_booth_integration_output_9_2), .A1 (
             nx8092), .S0 (nx35333)) ;
    mux21_ni ix8093 (.Y (nx8092), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_9_3), .S0 (nx36055)) ;
    mux21_ni ix18664 (.Y (nx18663), .A0 (booth_booth_integration_output_9_3), .A1 (
             nx8080), .S0 (nx35333)) ;
    mux21_ni ix8081 (.Y (nx8080), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_9_4), .S0 (nx36055)) ;
    mux21_ni ix18654 (.Y (nx18653), .A0 (booth_booth_integration_output_9_4), .A1 (
             nx8068), .S0 (nx35333)) ;
    mux21_ni ix8069 (.Y (nx8068), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_9_5), .S0 (nx36055)) ;
    mux21_ni ix18644 (.Y (nx18643), .A0 (booth_booth_integration_output_9_5), .A1 (
             nx8056), .S0 (nx35333)) ;
    mux21_ni ix8057 (.Y (nx8056), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_9_6), .S0 (nx36057)) ;
    mux21_ni ix18634 (.Y (nx18633), .A0 (booth_booth_integration_output_9_6), .A1 (
             nx8044), .S0 (nx35333)) ;
    mux21_ni ix8045 (.Y (nx8044), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_9_7), .S0 (nx36057)) ;
    mux21_ni ix18624 (.Y (nx18623), .A0 (booth_booth_integration_output_9_7), .A1 (
             nx8032), .S0 (nx36047)) ;
    mux21_ni ix8033 (.Y (nx8032), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_9_8), .S0 (nx36057)) ;
    mux21_ni ix18614 (.Y (nx18613), .A0 (booth_booth_integration_output_9_8), .A1 (
             nx8020), .S0 (nx36047)) ;
    mux21_ni ix8021 (.Y (nx8020), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_9_9), .S0 (nx36057)) ;
    mux21_ni ix18604 (.Y (nx18603), .A0 (booth_booth_integration_output_9_9), .A1 (
             nx8008), .S0 (nx36047)) ;
    mux21_ni ix8009 (.Y (nx8008), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_9_10), .S0 (nx36057)) ;
    mux21_ni ix18594 (.Y (nx18593), .A0 (booth_booth_integration_output_9_10), .A1 (
             nx7996), .S0 (nx36049)) ;
    mux21_ni ix7997 (.Y (nx7996), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_9_11), .S0 (nx36057)) ;
    mux21_ni ix18584 (.Y (nx18583), .A0 (booth_booth_integration_output_9_11), .A1 (
             nx7984), .S0 (nx36049)) ;
    mux21_ni ix7985 (.Y (nx7984), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_9_12), .S0 (nx36057)) ;
    mux21_ni ix18574 (.Y (nx18573), .A0 (booth_booth_integration_output_9_12), .A1 (
             nx7972), .S0 (nx36049)) ;
    mux21_ni ix7973 (.Y (nx7972), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_9_13), .S0 (nx36059)) ;
    mux21_ni ix18564 (.Y (nx18563), .A0 (booth_booth_integration_output_9_13), .A1 (
             nx7960), .S0 (nx36049)) ;
    mux21_ni ix7961 (.Y (nx7960), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_9_14), .S0 (nx36059)) ;
    mux21_ni ix18554 (.Y (nx18553), .A0 (booth_booth_integration_output_9_14), .A1 (
             nx7948), .S0 (nx36049)) ;
    mux21_ni ix7949 (.Y (nx7948), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_9_15), .S0 (nx36059)) ;
    mux21 ix18544 (.Y (nx18543), .A0 (nx27552), .A1 (nx27194), .S0 (nx36049)) ;
    mux21_ni ix18194 (.Y (nx18193), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_0), .A1 (nx34879), .S0 (
             nx35811)) ;
    and02 ix18180 (.Y (nx18179), .A0 (nx36345), .A1 (
          booth_booth_integrtaion_9_shift_Reg_count_0)) ;
    mux21_ni ix18374 (.Y (nx18373), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_9), .A1 (nx34865), .S0 (
             nx35811)) ;
    mux21_ni ix18364 (.Y (nx18363), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_8), .S0 (nx36049)) ;
    mux21_ni ix18354 (.Y (nx18353), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_8), .S0 (nx35811)) ;
    mux21_ni ix18344 (.Y (nx18343), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_7), .S0 (nx36051)) ;
    mux21_ni ix18334 (.Y (nx18333), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_7), .S0 (nx35811)) ;
    mux21_ni ix18324 (.Y (nx18323), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_6), .S0 (nx36051)) ;
    mux21_ni ix18314 (.Y (nx18313), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_6), .S0 (nx35811)) ;
    mux21_ni ix18304 (.Y (nx18303), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_5), .S0 (nx36051)) ;
    mux21_ni ix18294 (.Y (nx18293), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_5), .S0 (nx35811)) ;
    mux21_ni ix18284 (.Y (nx18283), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_4), .S0 (nx36051)) ;
    mux21_ni ix18274 (.Y (nx18273), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_4), .S0 (nx35813)) ;
    mux21_ni ix18264 (.Y (nx18263), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_3), .S0 (nx36051)) ;
    mux21_ni ix18254 (.Y (nx18253), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_3), .S0 (nx35813)) ;
    mux21_ni ix18244 (.Y (nx18243), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_2), .S0 (nx36051)) ;
    mux21_ni ix18234 (.Y (nx18233), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_2), .S0 (nx35813)) ;
    mux21_ni ix18224 (.Y (nx18223), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_1), .S0 (nx36051)) ;
    mux21_ni ix18214 (.Y (nx18213), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_9_shift_Reg_output_1), .S0 (nx35813)) ;
    mux21_ni ix18204 (.Y (nx18203), .A0 (
             booth_booth_integrtaion_9_shift_Reg_count_1), .A1 (nx34879), .S0 (
             nx36053)) ;
    and02 ix7389 (.Y (nx7388), .A0 (nx27267), .A1 (nx35759)) ;
    or03 ix27270 (.Y (nx27269), .A0 (nx27271), .A1 (
         booth_booth_integrtaion_9_shift_reg_output_0), .A2 (nx36345)) ;
    mux21_ni ix18534 (.Y (nx18533), .A0 (
             booth_booth_integrtaion_9_booth_output_16), .A1 (nx7918), .S0 (
             nx36053)) ;
    nor02ii ix7919 (.Y (nx7918), .A0 (nx27278), .A1 (nx36059)) ;
    nor02ii ix7395 (.Y (nx7394), .A0 (nx27262), .A1 (
            booth_booth_integrtaion_9_booth_output_16)) ;
    xor2 ix7913 (.Y (nx13149), .A0 (nx27284), .A1 (nx27548)) ;
    xor2 ix7901 (.Y (nx13151), .A0 (nx27309), .A1 (nx35339)) ;
    mux21_ni ix18514 (.Y (nx18513), .A0 (
             booth_booth_integrtaion_9_booth_output_18), .A1 (nx7894), .S0 (
             nx36053)) ;
    nor02ii ix7895 (.Y (nx7894), .A0 (nx27299), .A1 (nx36059)) ;
    xor2 ix7889 (.Y (nx13153), .A0 (nx27314), .A1 (nx27545)) ;
    or02 ix27331 (.Y (nx27330), .A0 (nx27267), .A1 (nx35761)) ;
    xor2 ix7877 (.Y (nx13155), .A0 (nx27348), .A1 (nx35341)) ;
    mux21_ni ix18494 (.Y (nx18493), .A0 (
             booth_booth_integrtaion_9_booth_output_20), .A1 (nx7870), .S0 (
             nx36053)) ;
    nor02ii ix7871 (.Y (nx7870), .A0 (nx27336), .A1 (nx36059)) ;
    xor2 ix7865 (.Y (nx13157), .A0 (nx27353), .A1 (nx27542)) ;
    xor2 ix7853 (.Y (nx13159), .A0 (nx27383), .A1 (nx35343)) ;
    mux21_ni ix18474 (.Y (nx18473), .A0 (
             booth_booth_integrtaion_9_booth_output_22), .A1 (nx7846), .S0 (
             nx36053)) ;
    nor02ii ix7847 (.Y (nx7846), .A0 (nx27371), .A1 (nx36059)) ;
    xor2 ix7841 (.Y (nx13161), .A0 (nx27388), .A1 (nx27539)) ;
    xor2 ix7829 (.Y (nx13162), .A0 (nx27418), .A1 (nx35345)) ;
    mux21_ni ix18454 (.Y (nx18453), .A0 (
             booth_booth_integrtaion_9_booth_output_24), .A1 (nx7822), .S0 (
             nx36053)) ;
    nor02ii ix7823 (.Y (nx7822), .A0 (nx27406), .A1 (nx36061)) ;
    xor2 ix7817 (.Y (nx13163), .A0 (nx27423), .A1 (nx27536)) ;
    xor2 ix7805 (.Y (nx13165), .A0 (nx27453), .A1 (nx35347)) ;
    mux21_ni ix18434 (.Y (nx18433), .A0 (
             booth_booth_integrtaion_9_booth_output_26), .A1 (nx7798), .S0 (
             nx36053)) ;
    nor02ii ix7799 (.Y (nx7798), .A0 (nx27441), .A1 (nx36061)) ;
    xor2 ix7793 (.Y (nx13167), .A0 (nx27458), .A1 (nx27533)) ;
    xor2 ix7781 (.Y (nx13169), .A0 (nx27488), .A1 (nx35349)) ;
    mux21_ni ix18414 (.Y (nx18413), .A0 (
             booth_booth_integrtaion_9_booth_output_28), .A1 (nx7774), .S0 (
             nx35331)) ;
    nor02ii ix7775 (.Y (nx7774), .A0 (nx27476), .A1 (nx36061)) ;
    xor2 ix7769 (.Y (nx13170), .A0 (nx27493), .A1 (nx27530)) ;
    xor2 ix7757 (.Y (nx13171), .A0 (nx27523), .A1 (nx35351)) ;
    mux21_ni ix18394 (.Y (nx18393), .A0 (
             booth_booth_integrtaion_9_booth_output_31), .A1 (nx7750), .S0 (
             nx35331)) ;
    nor02ii ix7751 (.Y (nx7750), .A0 (nx27511), .A1 (nx36061)) ;
    xor2 ix7745 (.Y (nx7744), .A0 (nx27523), .A1 (nx27526)) ;
    nor02ii ix7931 (.Y (nx7930), .A0 (nx7394), .A1 (nx36061)) ;
    or03 ix27577 (.Y (nx27576), .A0 (nx27760), .A1 (nx35843), .A2 (nx35361)) ;
    mux21_ni ix18984 (.Y (nx18983), .A0 (label_10_output[14]), .A1 (
             label_10_input_14), .S0 (nx36241)) ;
    mux21_ni ix8575 (.Y (nx8574), .A0 (nx8570), .A1 (
             label_10_input_state_machine_14), .S0 (nx35919)) ;
    mux21_ni ix18164 (.Y (nx18163), .A0 (label_10_input_state_machine_14), .A1 (
             mdr_data_out[158]), .S0 (nx36201)) ;
    mux21_ni ix18974 (.Y (nx18973), .A0 (label_10_output[13]), .A1 (
             label_10_input_13), .S0 (nx36241)) ;
    mux21_ni ix8549 (.Y (nx8548), .A0 (nx8544), .A1 (
             label_10_input_state_machine_13), .S0 (nx35921)) ;
    mux21_ni ix18964 (.Y (nx18963), .A0 (label_10_input_state_machine_13), .A1 (
             mdr_data_out[157]), .S0 (nx36201)) ;
    mux21_ni ix18934 (.Y (nx18933), .A0 (label_10_output[11]), .A1 (
             label_10_input_11), .S0 (nx36241)) ;
    mux21_ni ix8485 (.Y (nx8484), .A0 (nx8480), .A1 (
             label_10_input_state_machine_11), .S0 (nx35921)) ;
    mux21_ni ix18924 (.Y (nx18923), .A0 (label_10_input_state_machine_11), .A1 (
             mdr_data_out[155]), .S0 (nx36203)) ;
    mux21_ni ix18894 (.Y (nx18893), .A0 (label_10_output[9]), .A1 (
             label_10_input_9), .S0 (nx36241)) ;
    mux21_ni ix8421 (.Y (nx8420), .A0 (nx8416), .A1 (
             label_10_input_state_machine_9), .S0 (nx35921)) ;
    mux21_ni ix18884 (.Y (nx18883), .A0 (label_10_input_state_machine_9), .A1 (
             mdr_data_out[153]), .S0 (nx36203)) ;
    mux21_ni ix18854 (.Y (nx18853), .A0 (label_10_output[7]), .A1 (
             label_10_input_7), .S0 (nx36243)) ;
    mux21_ni ix8357 (.Y (nx8356), .A0 (nx8352), .A1 (
             label_10_input_state_machine_7), .S0 (nx35921)) ;
    mux21_ni ix18844 (.Y (nx18843), .A0 (label_10_input_state_machine_7), .A1 (
             mdr_data_out[151]), .S0 (nx36203)) ;
    mux21_ni ix18814 (.Y (nx18813), .A0 (label_10_output[5]), .A1 (
             label_10_input_5), .S0 (nx36243)) ;
    mux21_ni ix8293 (.Y (nx8292), .A0 (nx8288), .A1 (
             label_10_input_state_machine_5), .S0 (nx35921)) ;
    mux21_ni ix18804 (.Y (nx18803), .A0 (label_10_input_state_machine_5), .A1 (
             mdr_data_out[149]), .S0 (nx36203)) ;
    mux21_ni ix18774 (.Y (nx18773), .A0 (label_10_output[3]), .A1 (
             label_10_input_3), .S0 (nx36243)) ;
    mux21_ni ix8229 (.Y (nx8228), .A0 (nx8224), .A1 (
             label_10_input_state_machine_3), .S0 (nx35921)) ;
    mux21_ni ix18764 (.Y (nx18763), .A0 (label_10_input_state_machine_3), .A1 (
             mdr_data_out[147]), .S0 (nx36203)) ;
    mux21_ni ix18734 (.Y (nx18733), .A0 (label_10_output[1]), .A1 (
             label_10_input_1), .S0 (nx36243)) ;
    mux21_ni ix8165 (.Y (nx8164), .A0 (nx8160), .A1 (
             label_10_input_state_machine_1), .S0 (nx35921)) ;
    mux21_ni ix18724 (.Y (nx18723), .A0 (label_10_input_state_machine_1), .A1 (
             mdr_data_out[145]), .S0 (nx36203)) ;
    xnor2 ix27669 (.Y (nx27668), .A0 (nx27566), .A1 (nx27678)) ;
    mux21_ni ix18754 (.Y (nx18753), .A0 (label_10_output[2]), .A1 (
             label_10_input_2), .S0 (nx36243)) ;
    mux21_ni ix8197 (.Y (nx8196), .A0 (nx8192), .A1 (
             label_10_input_state_machine_2), .S0 (nx35923)) ;
    mux21_ni ix18744 (.Y (nx18743), .A0 (label_10_input_state_machine_2), .A1 (
             mdr_data_out[146]), .S0 (nx36203)) ;
    xnor2 ix27684 (.Y (nx27683), .A0 (nx27564), .A1 (nx27693)) ;
    mux21_ni ix18794 (.Y (nx18793), .A0 (label_10_output[4]), .A1 (
             label_10_input_4), .S0 (nx36243)) ;
    mux21_ni ix8261 (.Y (nx8260), .A0 (nx8256), .A1 (
             label_10_input_state_machine_4), .S0 (nx35923)) ;
    mux21_ni ix18784 (.Y (nx18783), .A0 (label_10_input_state_machine_4), .A1 (
             mdr_data_out[148]), .S0 (nx36205)) ;
    xnor2 ix27699 (.Y (nx27698), .A0 (nx27562), .A1 (nx27708)) ;
    mux21_ni ix18834 (.Y (nx18833), .A0 (label_10_output[6]), .A1 (
             label_10_input_6), .S0 (nx36243)) ;
    mux21_ni ix8325 (.Y (nx8324), .A0 (nx8320), .A1 (
             label_10_input_state_machine_6), .S0 (nx35923)) ;
    mux21_ni ix18824 (.Y (nx18823), .A0 (label_10_input_state_machine_6), .A1 (
             mdr_data_out[150]), .S0 (nx36205)) ;
    xnor2 ix27714 (.Y (nx27713), .A0 (nx27560), .A1 (nx27723)) ;
    mux21_ni ix18874 (.Y (nx18873), .A0 (label_10_output[8]), .A1 (
             label_10_input_8), .S0 (nx36245)) ;
    mux21_ni ix8389 (.Y (nx8388), .A0 (nx8384), .A1 (
             label_10_input_state_machine_8), .S0 (nx35923)) ;
    mux21_ni ix18864 (.Y (nx18863), .A0 (label_10_input_state_machine_8), .A1 (
             mdr_data_out[152]), .S0 (nx36205)) ;
    xnor2 ix27729 (.Y (nx27728), .A0 (nx27558), .A1 (nx27738)) ;
    mux21_ni ix18914 (.Y (nx18913), .A0 (label_10_output[10]), .A1 (
             label_10_input_10), .S0 (nx36245)) ;
    mux21_ni ix8453 (.Y (nx8452), .A0 (nx8448), .A1 (
             label_10_input_state_machine_10), .S0 (nx35923)) ;
    mux21_ni ix18904 (.Y (nx18903), .A0 (label_10_input_state_machine_10), .A1 (
             mdr_data_out[154]), .S0 (nx36205)) ;
    xnor2 ix27744 (.Y (nx27743), .A0 (nx27556), .A1 (nx27753)) ;
    mux21_ni ix18954 (.Y (nx18953), .A0 (label_10_output[12]), .A1 (
             label_10_input_12), .S0 (nx36245)) ;
    mux21_ni ix8517 (.Y (nx8516), .A0 (nx8512), .A1 (
             label_10_input_state_machine_12), .S0 (nx35923)) ;
    mux21_ni ix18944 (.Y (nx18943), .A0 (label_10_input_state_machine_12), .A1 (
             mdr_data_out[156]), .S0 (nx36205)) ;
    xnor2 ix27759 (.Y (nx27758), .A0 (nx27554), .A1 (nx27760)) ;
    or03 ix27766 (.Y (nx27765), .A0 (nx27949), .A1 (nx35843), .A2 (nx35361)) ;
    mux21_ni ix19274 (.Y (nx19273), .A0 (label_9_output[14]), .A1 (
             label_9_input_14), .S0 (nx36245)) ;
    mux21_ni ix9025 (.Y (nx9024), .A0 (nx9020), .A1 (
             label_9_input_state_machine_14), .S0 (nx35925)) ;
    mux21_ni ix19004 (.Y (nx19003), .A0 (label_9_input_state_machine_14), .A1 (
             mdr_data_out[142]), .S0 (nx36205)) ;
    mux21_ni ix19264 (.Y (nx19263), .A0 (label_9_output[13]), .A1 (
             label_9_input_13), .S0 (nx36245)) ;
    mux21_ni ix8999 (.Y (nx8998), .A0 (nx8994), .A1 (
             label_9_input_state_machine_13), .S0 (nx35925)) ;
    mux21_ni ix19254 (.Y (nx19253), .A0 (label_9_input_state_machine_13), .A1 (
             mdr_data_out[141]), .S0 (nx36205)) ;
    mux21_ni ix19224 (.Y (nx19223), .A0 (label_9_output[11]), .A1 (
             label_9_input_11), .S0 (nx36245)) ;
    mux21_ni ix8935 (.Y (nx8934), .A0 (nx8930), .A1 (
             label_9_input_state_machine_11), .S0 (nx35925)) ;
    mux21_ni ix19214 (.Y (nx19213), .A0 (label_9_input_state_machine_11), .A1 (
             mdr_data_out[139]), .S0 (nx36207)) ;
    mux21_ni ix19184 (.Y (nx19183), .A0 (label_9_output[9]), .A1 (
             label_9_input_9), .S0 (nx36245)) ;
    mux21_ni ix8871 (.Y (nx8870), .A0 (nx8866), .A1 (
             label_9_input_state_machine_9), .S0 (nx35925)) ;
    mux21_ni ix19174 (.Y (nx19173), .A0 (label_9_input_state_machine_9), .A1 (
             mdr_data_out[137]), .S0 (nx36207)) ;
    mux21_ni ix19144 (.Y (nx19143), .A0 (label_9_output[7]), .A1 (
             label_9_input_7), .S0 (nx36247)) ;
    mux21_ni ix8807 (.Y (nx8806), .A0 (nx8802), .A1 (
             label_9_input_state_machine_7), .S0 (nx35923)) ;
    mux21_ni ix19134 (.Y (nx19133), .A0 (label_9_input_state_machine_7), .A1 (
             mdr_data_out[135]), .S0 (nx36207)) ;
    mux21_ni ix19104 (.Y (nx19103), .A0 (label_9_output[5]), .A1 (
             label_9_input_5), .S0 (nx36247)) ;
    mux21_ni ix8743 (.Y (nx8742), .A0 (nx8738), .A1 (
             label_9_input_state_machine_5), .S0 (nx35165)) ;
    mux21_ni ix19094 (.Y (nx19093), .A0 (label_9_input_state_machine_5), .A1 (
             mdr_data_out[133]), .S0 (nx36207)) ;
    mux21_ni ix19064 (.Y (nx19063), .A0 (label_9_output[3]), .A1 (
             label_9_input_3), .S0 (nx36247)) ;
    mux21_ni ix8679 (.Y (nx8678), .A0 (nx8674), .A1 (
             label_9_input_state_machine_3), .S0 (nx35165)) ;
    mux21_ni ix19054 (.Y (nx19053), .A0 (label_9_input_state_machine_3), .A1 (
             mdr_data_out[131]), .S0 (nx36207)) ;
    mux21_ni ix19024 (.Y (nx19023), .A0 (label_9_output[1]), .A1 (
             label_9_input_1), .S0 (nx36247)) ;
    mux21_ni ix8615 (.Y (nx8614), .A0 (nx8610), .A1 (
             label_9_input_state_machine_1), .S0 (nx35165)) ;
    mux21_ni ix19014 (.Y (nx19013), .A0 (label_9_input_state_machine_1), .A1 (
             mdr_data_out[129]), .S0 (nx36207)) ;
    xnor2 ix27858 (.Y (nx27857), .A0 (nx27127), .A1 (nx27867)) ;
    mux21_ni ix19044 (.Y (nx19043), .A0 (label_9_output[2]), .A1 (
             label_9_input_2), .S0 (nx36247)) ;
    mux21_ni ix8647 (.Y (nx8646), .A0 (nx8642), .A1 (
             label_9_input_state_machine_2), .S0 (nx35165)) ;
    mux21_ni ix19034 (.Y (nx19033), .A0 (label_9_input_state_machine_2), .A1 (
             mdr_data_out[130]), .S0 (nx36207)) ;
    xnor2 ix27873 (.Y (nx27872), .A0 (nx27125), .A1 (nx27882)) ;
    mux21_ni ix19084 (.Y (nx19083), .A0 (label_9_output[4]), .A1 (
             label_9_input_4), .S0 (nx36247)) ;
    mux21_ni ix8711 (.Y (nx8710), .A0 (nx8706), .A1 (
             label_9_input_state_machine_4), .S0 (nx35165)) ;
    mux21_ni ix19074 (.Y (nx19073), .A0 (label_9_input_state_machine_4), .A1 (
             mdr_data_out[132]), .S0 (nx36209)) ;
    xnor2 ix27888 (.Y (nx27887), .A0 (nx27123), .A1 (nx27897)) ;
    mux21_ni ix19124 (.Y (nx19123), .A0 (label_9_output[6]), .A1 (
             label_9_input_6), .S0 (nx36247)) ;
    mux21_ni ix8775 (.Y (nx8774), .A0 (nx8770), .A1 (
             label_9_input_state_machine_6), .S0 (nx35165)) ;
    mux21_ni ix19114 (.Y (nx19113), .A0 (label_9_input_state_machine_6), .A1 (
             mdr_data_out[134]), .S0 (nx36209)) ;
    xnor2 ix27903 (.Y (nx27902), .A0 (nx27121), .A1 (nx27912)) ;
    mux21_ni ix19164 (.Y (nx19163), .A0 (label_9_output[8]), .A1 (
             label_9_input_8), .S0 (nx36249)) ;
    mux21_ni ix8839 (.Y (nx8838), .A0 (nx8834), .A1 (
             label_9_input_state_machine_8), .S0 (nx35165)) ;
    mux21_ni ix19154 (.Y (nx19153), .A0 (label_9_input_state_machine_8), .A1 (
             mdr_data_out[136]), .S0 (nx36209)) ;
    xnor2 ix27918 (.Y (nx27917), .A0 (nx27119), .A1 (nx27927)) ;
    mux21_ni ix19204 (.Y (nx19203), .A0 (label_9_output[10]), .A1 (
             label_9_input_10), .S0 (nx36249)) ;
    mux21_ni ix8903 (.Y (nx8902), .A0 (nx8898), .A1 (
             label_9_input_state_machine_10), .S0 (nx35925)) ;
    mux21_ni ix19194 (.Y (nx19193), .A0 (label_9_input_state_machine_10), .A1 (
             mdr_data_out[138]), .S0 (nx36209)) ;
    xnor2 ix27933 (.Y (nx27932), .A0 (nx27117), .A1 (nx27942)) ;
    mux21_ni ix19244 (.Y (nx19243), .A0 (label_9_output[12]), .A1 (
             label_9_input_12), .S0 (nx36249)) ;
    mux21_ni ix8967 (.Y (nx8966), .A0 (nx8962), .A1 (
             label_9_input_state_machine_12), .S0 (nx35927)) ;
    mux21_ni ix19234 (.Y (nx19233), .A0 (label_9_input_state_machine_12), .A1 (
             mdr_data_out[140]), .S0 (nx36209)) ;
    xnor2 ix27948 (.Y (nx27947), .A0 (nx27115), .A1 (nx27949)) ;
    xnor2 ix9045 (.Y (nx9044), .A0 (nx27573), .A1 (nx27763)) ;
    xnor2 ix27953 (.Y (nx27952), .A0 (nx27956), .A1 (
          max_calc_comparator_fifth_inp1_13)) ;
    or03 ix27971 (.Y (nx27970), .A0 (nx27753), .A1 (nx35845), .A2 (nx35361)) ;
    or03 ix27977 (.Y (nx27976), .A0 (nx27942), .A1 (nx35845), .A2 (nx35361)) ;
    xnor2 ix9081 (.Y (nx9080), .A0 (nx27967), .A1 (nx27974)) ;
    xnor2 ix27981 (.Y (nx27980), .A0 (nx27984), .A1 (
          max_calc_comparator_fifth_inp1_11)) ;
    or03 ix27999 (.Y (nx27998), .A0 (nx27738), .A1 (nx35845), .A2 (nx36065)) ;
    or03 ix28005 (.Y (nx28004), .A0 (nx27927), .A1 (nx35845), .A2 (nx36065)) ;
    xnor2 ix9117 (.Y (nx9116), .A0 (nx27995), .A1 (nx28002)) ;
    xnor2 ix28009 (.Y (nx28008), .A0 (nx28012), .A1 (
          max_calc_comparator_fifth_inp1_9)) ;
    or03 ix28027 (.Y (nx28026), .A0 (nx27723), .A1 (nx35845), .A2 (nx36065)) ;
    or03 ix28033 (.Y (nx28032), .A0 (nx27912), .A1 (nx35845), .A2 (nx36065)) ;
    xnor2 ix9153 (.Y (nx9152), .A0 (nx28023), .A1 (nx28030)) ;
    xnor2 ix28037 (.Y (nx28036), .A0 (nx28040), .A1 (
          max_calc_comparator_fifth_inp1_7)) ;
    or03 ix28055 (.Y (nx28054), .A0 (nx27708), .A1 (nx35845), .A2 (nx36065)) ;
    or03 ix28061 (.Y (nx28060), .A0 (nx27897), .A1 (nx35847), .A2 (nx36065)) ;
    xnor2 ix9189 (.Y (nx9188), .A0 (nx28051), .A1 (nx28058)) ;
    xnor2 ix28065 (.Y (nx28064), .A0 (nx28068), .A1 (
          max_calc_comparator_fifth_inp1_5)) ;
    or03 ix28083 (.Y (nx28082), .A0 (nx27693), .A1 (nx35847), .A2 (nx36065)) ;
    or03 ix28089 (.Y (nx28088), .A0 (nx27882), .A1 (nx35847), .A2 (nx35363)) ;
    xnor2 ix9225 (.Y (nx9224), .A0 (nx28079), .A1 (nx28086)) ;
    xnor2 ix28093 (.Y (nx28092), .A0 (nx28096), .A1 (
          max_calc_comparator_fifth_inp1_3)) ;
    or03 ix28111 (.Y (nx28110), .A0 (nx27678), .A1 (nx35847), .A2 (nx35363)) ;
    or03 ix28117 (.Y (nx28116), .A0 (nx27867), .A1 (nx35847), .A2 (nx35363)) ;
    xnor2 ix9261 (.Y (nx9260), .A0 (nx28107), .A1 (nx28114)) ;
    xnor2 ix9279 (.Y (nx9278), .A0 (nx28122), .A1 (nx28126)) ;
    xnor2 ix9489 (.Y (nx9488), .A0 (nx28137), .A1 (nx28155)) ;
    mux21_ni ix19574 (.Y (nx19573), .A0 (label_10_output[15]), .A1 (
             label_10_input_15), .S0 (nx36249)) ;
    mux21_ni ix9429 (.Y (nx9428), .A0 (nx9424), .A1 (
             label_10_input_state_machine_15), .S0 (nx35927)) ;
    mux21_ni ix19564 (.Y (nx19563), .A0 (label_10_input_state_machine_15), .A1 (
             mdr_data_out[159]), .S0 (nx36209)) ;
    xor2 ix28151 (.Y (nx28150), .A0 (nx27552), .A1 (label_10_output[15])) ;
    mux21_ni ix19604 (.Y (nx19603), .A0 (label_9_output[15]), .A1 (
             label_9_input_15), .S0 (nx36249)) ;
    mux21_ni ix9469 (.Y (nx9468), .A0 (nx9464), .A1 (
             label_9_input_state_machine_15), .S0 (nx35927)) ;
    mux21_ni ix19594 (.Y (nx19593), .A0 (label_9_input_state_machine_15), .A1 (
             mdr_data_out[143]), .S0 (nx36209)) ;
    xor2 ix28169 (.Y (nx28168), .A0 (nx27113), .A1 (label_9_output[15])) ;
    or04 ix28173 (.Y (nx28172), .A0 (rst), .A1 (nx26180), .A2 (max_calc_state_3)
         , .A3 (nx26188)) ;
    mux21_ni ix25474 (.Y (nx25473), .A0 (max_calc_comparator_first_inp2_0), .A1 (
             nx18892), .S0 (nx36281)) ;
    mux21_ni ix18893 (.Y (nx18892), .A0 (nx18888), .A1 (nx18864), .S0 (nx35965)
             ) ;
    mux21_ni ix18865 (.Y (nx18864), .A0 (max_calc_ans2_0), .A1 (
             label_2_output[0]), .S0 (nx35987)) ;
    mux21_ni ix16374 (.Y (nx16373), .A0 (label_2_output[0]), .A1 (
             label_2_input_0), .S0 (nx36249)) ;
    mux21_ni ix16364 (.Y (nx16363), .A0 (label_2_input_state_machine_0), .A1 (
             mdr_data_out[16]), .S0 (nx36211)) ;
    mux21_ni ix16354 (.Y (nx16353), .A0 (nx35727), .A1 (nx4398), .S0 (nx35379)
             ) ;
    mux21_ni ix4399 (.Y (nx4398), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_1_1), .S0 (nx36085)) ;
    mux21_ni ix16344 (.Y (nx16343), .A0 (booth_booth_integration_output_1_1), .A1 (
             nx4386), .S0 (nx35379)) ;
    mux21_ni ix4387 (.Y (nx4386), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_1_2), .S0 (nx36085)) ;
    mux21_ni ix16334 (.Y (nx16333), .A0 (booth_booth_integration_output_1_2), .A1 (
             nx4374), .S0 (nx35379)) ;
    mux21_ni ix4375 (.Y (nx4374), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_1_3), .S0 (nx36085)) ;
    mux21_ni ix16324 (.Y (nx16323), .A0 (booth_booth_integration_output_1_3), .A1 (
             nx4362), .S0 (nx35379)) ;
    mux21_ni ix4363 (.Y (nx4362), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_1_4), .S0 (nx36085)) ;
    mux21_ni ix16314 (.Y (nx16313), .A0 (booth_booth_integration_output_1_4), .A1 (
             nx4350), .S0 (nx35379)) ;
    mux21_ni ix4351 (.Y (nx4350), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_1_5), .S0 (nx36085)) ;
    mux21_ni ix16304 (.Y (nx16303), .A0 (booth_booth_integration_output_1_5), .A1 (
             nx4338), .S0 (nx35379)) ;
    mux21_ni ix4339 (.Y (nx4338), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_1_6), .S0 (nx36087)) ;
    mux21_ni ix16294 (.Y (nx16293), .A0 (booth_booth_integration_output_1_6), .A1 (
             nx4326), .S0 (nx35379)) ;
    mux21_ni ix4327 (.Y (nx4326), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_1_7), .S0 (nx36087)) ;
    mux21_ni ix16284 (.Y (nx16283), .A0 (booth_booth_integration_output_1_7), .A1 (
             nx4314), .S0 (nx36077)) ;
    mux21_ni ix4315 (.Y (nx4314), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_1_8), .S0 (nx36087)) ;
    mux21_ni ix16274 (.Y (nx16273), .A0 (booth_booth_integration_output_1_8), .A1 (
             nx4302), .S0 (nx36077)) ;
    mux21_ni ix4303 (.Y (nx4302), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_1_9), .S0 (nx36087)) ;
    mux21_ni ix16264 (.Y (nx16263), .A0 (booth_booth_integration_output_1_9), .A1 (
             nx4290), .S0 (nx36077)) ;
    mux21_ni ix4291 (.Y (nx4290), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_1_10), .S0 (nx36087)) ;
    mux21_ni ix16254 (.Y (nx16253), .A0 (booth_booth_integration_output_1_10), .A1 (
             nx4278), .S0 (nx36079)) ;
    mux21_ni ix4279 (.Y (nx4278), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_1_11), .S0 (nx36087)) ;
    mux21_ni ix16244 (.Y (nx16243), .A0 (booth_booth_integration_output_1_11), .A1 (
             nx4266), .S0 (nx36079)) ;
    mux21_ni ix4267 (.Y (nx4266), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_1_12), .S0 (nx36087)) ;
    mux21_ni ix16234 (.Y (nx16233), .A0 (booth_booth_integration_output_1_12), .A1 (
             nx4254), .S0 (nx36079)) ;
    mux21_ni ix4255 (.Y (nx4254), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_1_13), .S0 (nx36089)) ;
    mux21_ni ix16224 (.Y (nx16223), .A0 (booth_booth_integration_output_1_13), .A1 (
             nx4242), .S0 (nx36079)) ;
    mux21_ni ix4243 (.Y (nx4242), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_1_14), .S0 (nx36089)) ;
    mux21_ni ix16214 (.Y (nx16213), .A0 (booth_booth_integration_output_1_14), .A1 (
             nx4230), .S0 (nx36079)) ;
    mux21_ni ix4231 (.Y (nx4230), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_1_15), .S0 (nx36089)) ;
    mux21 ix16204 (.Y (nx16203), .A0 (nx28594), .A1 (nx28236), .S0 (nx36079)) ;
    mux21_ni ix15854 (.Y (nx15853), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_0), .A1 (nx34635), .S0 (
             nx35815)) ;
    and02 ix15840 (.Y (nx15839), .A0 (nx36323), .A1 (
          booth_booth_integrtaion_1_shift_Reg_count_0)) ;
    mux21_ni ix16034 (.Y (nx16033), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_9), .A1 (nx34621), .S0 (
             nx35815)) ;
    mux21_ni ix16024 (.Y (nx16023), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_8), .S0 (nx36079)) ;
    mux21_ni ix16014 (.Y (nx16013), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_8), .S0 (nx35815)) ;
    mux21_ni ix16004 (.Y (nx16003), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_7), .S0 (nx36081)) ;
    mux21_ni ix15994 (.Y (nx15993), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_7), .S0 (nx35815)) ;
    mux21_ni ix15984 (.Y (nx15983), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_6), .S0 (nx36081)) ;
    mux21_ni ix15974 (.Y (nx15973), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_6), .S0 (nx35815)) ;
    mux21_ni ix15964 (.Y (nx15963), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_5), .S0 (nx36081)) ;
    mux21_ni ix15954 (.Y (nx15953), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_5), .S0 (nx35815)) ;
    mux21_ni ix15944 (.Y (nx15943), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_4), .S0 (nx36081)) ;
    mux21_ni ix15934 (.Y (nx15933), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_4), .S0 (nx35817)) ;
    mux21_ni ix15924 (.Y (nx15923), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_3), .S0 (nx36081)) ;
    mux21_ni ix15914 (.Y (nx15913), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_3), .S0 (nx35817)) ;
    mux21_ni ix15904 (.Y (nx15903), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_2), .S0 (nx36081)) ;
    mux21_ni ix15894 (.Y (nx15893), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_2), .S0 (nx35817)) ;
    mux21_ni ix15884 (.Y (nx15883), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_1), .S0 (nx36081)) ;
    mux21_ni ix15874 (.Y (nx15873), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_1_shift_Reg_output_1), .S0 (nx35817)) ;
    mux21_ni ix15864 (.Y (nx15863), .A0 (
             booth_booth_integrtaion_1_shift_Reg_count_1), .A1 (nx34635), .S0 (
             nx36083)) ;
    and02 ix3671 (.Y (nx3670), .A0 (nx28309), .A1 (nx35727)) ;
    or03 ix28312 (.Y (nx28311), .A0 (nx28313), .A1 (
         booth_booth_integrtaion_1_shift_reg_output_0), .A2 (nx36323)) ;
    mux21_ni ix16194 (.Y (nx16193), .A0 (
             booth_booth_integrtaion_1_booth_output_16), .A1 (nx4200), .S0 (
             nx36083)) ;
    nor02ii ix4201 (.Y (nx4200), .A0 (nx28320), .A1 (nx36089)) ;
    nor02ii ix3677 (.Y (nx3676), .A0 (nx28304), .A1 (
            booth_booth_integrtaion_1_booth_output_16)) ;
    xor2 ix4195 (.Y (nx13017), .A0 (nx28326), .A1 (nx28590)) ;
    xor2 ix4183 (.Y (nx13018), .A0 (nx28351), .A1 (nx35385)) ;
    mux21_ni ix16174 (.Y (nx16173), .A0 (
             booth_booth_integrtaion_1_booth_output_18), .A1 (nx4176), .S0 (
             nx36083)) ;
    nor02ii ix4177 (.Y (nx4176), .A0 (nx28341), .A1 (nx36089)) ;
    xor2 ix4171 (.Y (nx13019), .A0 (nx28356), .A1 (nx28587)) ;
    or02 ix28373 (.Y (nx28372), .A0 (nx28309), .A1 (nx35729)) ;
    xor2 ix4159 (.Y (nx13021), .A0 (nx28390), .A1 (nx35387)) ;
    mux21_ni ix16154 (.Y (nx16153), .A0 (
             booth_booth_integrtaion_1_booth_output_20), .A1 (nx4152), .S0 (
             nx36083)) ;
    nor02ii ix4153 (.Y (nx4152), .A0 (nx28378), .A1 (nx36089)) ;
    xor2 ix4147 (.Y (nx13023), .A0 (nx28395), .A1 (nx28584)) ;
    xor2 ix4135 (.Y (nx13025), .A0 (nx28425), .A1 (nx35389)) ;
    mux21_ni ix16134 (.Y (nx16133), .A0 (
             booth_booth_integrtaion_1_booth_output_22), .A1 (nx4128), .S0 (
             nx36083)) ;
    nor02ii ix4129 (.Y (nx4128), .A0 (nx28413), .A1 (nx36089)) ;
    xor2 ix4123 (.Y (nx13026), .A0 (nx28430), .A1 (nx28581)) ;
    xor2 ix4111 (.Y (nx13027), .A0 (nx28460), .A1 (nx35391)) ;
    mux21_ni ix16114 (.Y (nx16113), .A0 (
             booth_booth_integrtaion_1_booth_output_24), .A1 (nx4104), .S0 (
             nx36083)) ;
    nor02ii ix4105 (.Y (nx4104), .A0 (nx28448), .A1 (nx36091)) ;
    xor2 ix4099 (.Y (nx13029), .A0 (nx28465), .A1 (nx28578)) ;
    xor2 ix4087 (.Y (nx13031), .A0 (nx28495), .A1 (nx35393)) ;
    mux21_ni ix16094 (.Y (nx16093), .A0 (
             booth_booth_integrtaion_1_booth_output_26), .A1 (nx4080), .S0 (
             nx36083)) ;
    nor02ii ix4081 (.Y (nx4080), .A0 (nx28483), .A1 (nx36091)) ;
    xor2 ix4075 (.Y (nx13033), .A0 (nx28500), .A1 (nx28575)) ;
    xor2 ix4063 (.Y (nx13035), .A0 (nx28530), .A1 (nx35395)) ;
    mux21_ni ix16074 (.Y (nx16073), .A0 (
             booth_booth_integrtaion_1_booth_output_28), .A1 (nx4056), .S0 (
             nx35377)) ;
    nor02ii ix4057 (.Y (nx4056), .A0 (nx28518), .A1 (nx36091)) ;
    xor2 ix4051 (.Y (nx13037), .A0 (nx28535), .A1 (nx28572)) ;
    xor2 ix4039 (.Y (nx13039), .A0 (nx28565), .A1 (nx35397)) ;
    mux21_ni ix16054 (.Y (nx16053), .A0 (
             booth_booth_integrtaion_1_booth_output_31), .A1 (nx4032), .S0 (
             nx35377)) ;
    nor02ii ix4033 (.Y (nx4032), .A0 (nx28553), .A1 (nx36091)) ;
    xor2 ix4027 (.Y (nx4026), .A0 (nx28565), .A1 (nx28568)) ;
    nor02ii ix4213 (.Y (nx4212), .A0 (nx3676), .A1 (nx36091)) ;
    mux21_ni ix25444 (.Y (nx25443), .A0 (nx18854), .A1 (max_calc_ans2_0), .S0 (
             nx35851)) ;
    mux21 ix18855 (.Y (nx18854), .A0 (nx30546), .A1 (nx28617), .S0 (nx35899)) ;
    mux21_ni ix16933 (.Y (nx16932), .A0 (max_calc_ans3_0), .A1 (
             label_3_output[0]), .S0 (nx35977)) ;
    mux21_ni ix15524 (.Y (nx15523), .A0 (label_3_output[0]), .A1 (
             label_3_input_0), .S0 (nx36249)) ;
    mux21_ni ix15514 (.Y (nx15513), .A0 (label_3_input_state_machine_0), .A1 (
             mdr_data_out[32]), .S0 (nx36211)) ;
    mux21_ni ix15504 (.Y (nx15503), .A0 (nx35723), .A1 (nx3060), .S0 (nx35405)
             ) ;
    mux21_ni ix3061 (.Y (nx3060), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_2_1), .S0 (nx36101)) ;
    mux21_ni ix15494 (.Y (nx15493), .A0 (booth_booth_integration_output_2_1), .A1 (
             nx3048), .S0 (nx35405)) ;
    mux21_ni ix3049 (.Y (nx3048), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_2_2), .S0 (nx36101)) ;
    mux21_ni ix15484 (.Y (nx15483), .A0 (booth_booth_integration_output_2_2), .A1 (
             nx3036), .S0 (nx35405)) ;
    mux21_ni ix3037 (.Y (nx3036), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_2_3), .S0 (nx36101)) ;
    mux21_ni ix15474 (.Y (nx15473), .A0 (booth_booth_integration_output_2_3), .A1 (
             nx3024), .S0 (nx35405)) ;
    mux21_ni ix3025 (.Y (nx3024), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_2_4), .S0 (nx36101)) ;
    mux21_ni ix15464 (.Y (nx15463), .A0 (booth_booth_integration_output_2_4), .A1 (
             nx3012), .S0 (nx35405)) ;
    mux21_ni ix3013 (.Y (nx3012), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_2_5), .S0 (nx36101)) ;
    mux21_ni ix15454 (.Y (nx15453), .A0 (booth_booth_integration_output_2_5), .A1 (
             nx3000), .S0 (nx35405)) ;
    mux21_ni ix3001 (.Y (nx3000), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_2_6), .S0 (nx36103)) ;
    mux21_ni ix15444 (.Y (nx15443), .A0 (booth_booth_integration_output_2_6), .A1 (
             nx2988), .S0 (nx35405)) ;
    mux21_ni ix2989 (.Y (nx2988), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_2_7), .S0 (nx36103)) ;
    mux21_ni ix15434 (.Y (nx15433), .A0 (booth_booth_integration_output_2_7), .A1 (
             nx2976), .S0 (nx36093)) ;
    mux21_ni ix2977 (.Y (nx2976), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_2_8), .S0 (nx36103)) ;
    mux21_ni ix15424 (.Y (nx15423), .A0 (booth_booth_integration_output_2_8), .A1 (
             nx2964), .S0 (nx36093)) ;
    mux21_ni ix2965 (.Y (nx2964), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_2_9), .S0 (nx36103)) ;
    mux21_ni ix15414 (.Y (nx15413), .A0 (booth_booth_integration_output_2_9), .A1 (
             nx2952), .S0 (nx36093)) ;
    mux21_ni ix2953 (.Y (nx2952), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_2_10), .S0 (nx36103)) ;
    mux21_ni ix15404 (.Y (nx15403), .A0 (booth_booth_integration_output_2_10), .A1 (
             nx2940), .S0 (nx36095)) ;
    mux21_ni ix2941 (.Y (nx2940), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_2_11), .S0 (nx36103)) ;
    mux21_ni ix15394 (.Y (nx15393), .A0 (booth_booth_integration_output_2_11), .A1 (
             nx2928), .S0 (nx36095)) ;
    mux21_ni ix2929 (.Y (nx2928), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_2_12), .S0 (nx36103)) ;
    mux21_ni ix15384 (.Y (nx15383), .A0 (booth_booth_integration_output_2_12), .A1 (
             nx2916), .S0 (nx36095)) ;
    mux21_ni ix2917 (.Y (nx2916), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_2_13), .S0 (nx36105)) ;
    mux21_ni ix15374 (.Y (nx15373), .A0 (booth_booth_integration_output_2_13), .A1 (
             nx2904), .S0 (nx36095)) ;
    mux21_ni ix2905 (.Y (nx2904), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_2_14), .S0 (nx36105)) ;
    mux21_ni ix15364 (.Y (nx15363), .A0 (booth_booth_integration_output_2_14), .A1 (
             nx2892), .S0 (nx36095)) ;
    mux21_ni ix2893 (.Y (nx2892), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_2_15), .S0 (nx36105)) ;
    mux21 ix15354 (.Y (nx15353), .A0 (nx29037), .A1 (nx28679), .S0 (nx36095)) ;
    mux21_ni ix15004 (.Y (nx15003), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_0), .A1 (nx34603), .S0 (
             nx35819)) ;
    and02 ix14990 (.Y (nx14989), .A0 (nx36319), .A1 (
          booth_booth_integrtaion_2_shift_Reg_count_0)) ;
    mux21_ni ix15184 (.Y (nx15183), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_9), .A1 (nx34589), .S0 (
             nx35819)) ;
    mux21_ni ix15174 (.Y (nx15173), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_8), .S0 (nx36095)) ;
    mux21_ni ix15164 (.Y (nx15163), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_8), .S0 (nx35819)) ;
    mux21_ni ix15154 (.Y (nx15153), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_7), .S0 (nx36097)) ;
    mux21_ni ix15144 (.Y (nx15143), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_7), .S0 (nx35819)) ;
    mux21_ni ix15134 (.Y (nx15133), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_6), .S0 (nx36097)) ;
    mux21_ni ix15124 (.Y (nx15123), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_6), .S0 (nx35819)) ;
    mux21_ni ix15114 (.Y (nx15113), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_5), .S0 (nx36097)) ;
    mux21_ni ix15104 (.Y (nx15103), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_5), .S0 (nx35819)) ;
    mux21_ni ix15094 (.Y (nx15093), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_4), .S0 (nx36097)) ;
    mux21_ni ix15084 (.Y (nx15083), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_4), .S0 (nx35821)) ;
    mux21_ni ix15074 (.Y (nx15073), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_3), .S0 (nx36097)) ;
    mux21_ni ix15064 (.Y (nx15063), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_3), .S0 (nx35821)) ;
    mux21_ni ix15054 (.Y (nx15053), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_2), .S0 (nx36097)) ;
    mux21_ni ix15044 (.Y (nx15043), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_2), .S0 (nx35821)) ;
    mux21_ni ix15034 (.Y (nx15033), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_1), .S0 (nx36097)) ;
    mux21_ni ix15024 (.Y (nx15023), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_2_shift_Reg_output_1), .S0 (nx35821)) ;
    mux21_ni ix15014 (.Y (nx15013), .A0 (
             booth_booth_integrtaion_2_shift_Reg_count_1), .A1 (nx34603), .S0 (
             nx36099)) ;
    and02 ix2333 (.Y (nx2332), .A0 (nx28752), .A1 (nx35723)) ;
    or03 ix28755 (.Y (nx28754), .A0 (nx28756), .A1 (
         booth_booth_integrtaion_2_shift_reg_output_0), .A2 (nx36319)) ;
    mux21_ni ix15344 (.Y (nx15343), .A0 (
             booth_booth_integrtaion_2_booth_output_16), .A1 (nx2862), .S0 (
             nx36099)) ;
    nor02ii ix2863 (.Y (nx2862), .A0 (nx28763), .A1 (nx36105)) ;
    nor02ii ix2339 (.Y (nx2338), .A0 (nx28747), .A1 (
            booth_booth_integrtaion_2_booth_output_16)) ;
    xor2 ix2857 (.Y (nx12965), .A0 (nx28769), .A1 (nx29033)) ;
    xor2 ix2845 (.Y (nx12967), .A0 (nx28794), .A1 (nx35411)) ;
    mux21_ni ix15324 (.Y (nx15323), .A0 (
             booth_booth_integrtaion_2_booth_output_18), .A1 (nx2838), .S0 (
             nx36099)) ;
    nor02ii ix2839 (.Y (nx2838), .A0 (nx28784), .A1 (nx36105)) ;
    xor2 ix2833 (.Y (nx12969), .A0 (nx28799), .A1 (nx29030)) ;
    or02 ix28816 (.Y (nx28815), .A0 (nx28752), .A1 (nx35725)) ;
    xor2 ix2821 (.Y (nx12970), .A0 (nx28833), .A1 (nx35413)) ;
    mux21_ni ix15304 (.Y (nx15303), .A0 (
             booth_booth_integrtaion_2_booth_output_20), .A1 (nx2814), .S0 (
             nx36099)) ;
    nor02ii ix2815 (.Y (nx2814), .A0 (nx28821), .A1 (nx36105)) ;
    xor2 ix2809 (.Y (nx12971), .A0 (nx28838), .A1 (nx29027)) ;
    xor2 ix2797 (.Y (nx12973), .A0 (nx28868), .A1 (nx35415)) ;
    mux21_ni ix15284 (.Y (nx15283), .A0 (
             booth_booth_integrtaion_2_booth_output_22), .A1 (nx2790), .S0 (
             nx36099)) ;
    nor02ii ix2791 (.Y (nx2790), .A0 (nx28856), .A1 (nx36105)) ;
    xor2 ix2785 (.Y (nx12975), .A0 (nx28873), .A1 (nx29024)) ;
    xor2 ix2773 (.Y (nx12977), .A0 (nx28903), .A1 (nx35417)) ;
    mux21_ni ix15264 (.Y (nx15263), .A0 (
             booth_booth_integrtaion_2_booth_output_24), .A1 (nx2766), .S0 (
             nx36099)) ;
    nor02ii ix2767 (.Y (nx2766), .A0 (nx28891), .A1 (nx36107)) ;
    xor2 ix2761 (.Y (nx12978), .A0 (nx28908), .A1 (nx29021)) ;
    xor2 ix2749 (.Y (nx12979), .A0 (nx28938), .A1 (nx35419)) ;
    mux21_ni ix15244 (.Y (nx15243), .A0 (
             booth_booth_integrtaion_2_booth_output_26), .A1 (nx2742), .S0 (
             nx36099)) ;
    nor02ii ix2743 (.Y (nx2742), .A0 (nx28926), .A1 (nx36107)) ;
    xor2 ix2737 (.Y (nx12981), .A0 (nx28943), .A1 (nx29018)) ;
    xor2 ix2725 (.Y (nx12983), .A0 (nx28973), .A1 (nx35421)) ;
    mux21_ni ix15224 (.Y (nx15223), .A0 (
             booth_booth_integrtaion_2_booth_output_28), .A1 (nx2718), .S0 (
             nx35403)) ;
    nor02ii ix2719 (.Y (nx2718), .A0 (nx28961), .A1 (nx36107)) ;
    xor2 ix2713 (.Y (nx12985), .A0 (nx28978), .A1 (nx29015)) ;
    xor2 ix2701 (.Y (nx12987), .A0 (nx29008), .A1 (nx35423)) ;
    mux21_ni ix15204 (.Y (nx15203), .A0 (
             booth_booth_integrtaion_2_booth_output_31), .A1 (nx2694), .S0 (
             nx35403)) ;
    nor02ii ix2695 (.Y (nx2694), .A0 (nx28996), .A1 (nx36107)) ;
    xor2 ix2689 (.Y (nx2688), .A0 (nx29008), .A1 (nx29011)) ;
    nor02ii ix2875 (.Y (nx2874), .A0 (nx2338), .A1 (nx36107)) ;
    ao32 ix24264 (.Y (nx24263), .A0 (nx35959), .A1 (nx35645), .A2 (nx36291), .B0 (
         max_calc_ans3_0), .B1 (nx35877)) ;
    mux21 ix29058 (.Y (nx35645), .A0 (nx29502), .A1 (nx29061), .S0 (nx35887)) ;
    mux21_ni ix20194 (.Y (nx20193), .A0 (label_5_output[0]), .A1 (
             label_5_input_0), .S0 (nx36251)) ;
    mux21_ni ix20184 (.Y (nx20183), .A0 (label_5_input_state_machine_0), .A1 (
             mdr_data_out[64]), .S0 (nx36211)) ;
    mux21_ni ix20174 (.Y (nx20173), .A0 (nx35763), .A1 (nx10374), .S0 (nx35431)
             ) ;
    mux21_ni ix10375 (.Y (nx10374), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_4_1), .S0 (nx36117)) ;
    mux21_ni ix20164 (.Y (nx20163), .A0 (booth_booth_integration_output_4_1), .A1 (
             nx10362), .S0 (nx35431)) ;
    mux21_ni ix10363 (.Y (nx10362), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_4_2), .S0 (nx36117)) ;
    mux21_ni ix20154 (.Y (nx20153), .A0 (booth_booth_integration_output_4_2), .A1 (
             nx10350), .S0 (nx35431)) ;
    mux21_ni ix10351 (.Y (nx10350), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_4_3), .S0 (nx36117)) ;
    mux21_ni ix20144 (.Y (nx20143), .A0 (booth_booth_integration_output_4_3), .A1 (
             nx10338), .S0 (nx35431)) ;
    mux21_ni ix10339 (.Y (nx10338), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_4_4), .S0 (nx36117)) ;
    mux21_ni ix20134 (.Y (nx20133), .A0 (booth_booth_integration_output_4_4), .A1 (
             nx10326), .S0 (nx35431)) ;
    mux21_ni ix10327 (.Y (nx10326), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_4_5), .S0 (nx36117)) ;
    mux21_ni ix20124 (.Y (nx20123), .A0 (booth_booth_integration_output_4_5), .A1 (
             nx10314), .S0 (nx35431)) ;
    mux21_ni ix10315 (.Y (nx10314), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_4_6), .S0 (nx36119)) ;
    mux21_ni ix20114 (.Y (nx20113), .A0 (booth_booth_integration_output_4_6), .A1 (
             nx10302), .S0 (nx35431)) ;
    mux21_ni ix10303 (.Y (nx10302), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_4_7), .S0 (nx36119)) ;
    mux21_ni ix20104 (.Y (nx20103), .A0 (booth_booth_integration_output_4_7), .A1 (
             nx10290), .S0 (nx36109)) ;
    mux21_ni ix10291 (.Y (nx10290), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_4_8), .S0 (nx36119)) ;
    mux21_ni ix20094 (.Y (nx20093), .A0 (booth_booth_integration_output_4_8), .A1 (
             nx10278), .S0 (nx36109)) ;
    mux21_ni ix10279 (.Y (nx10278), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_4_9), .S0 (nx36119)) ;
    mux21_ni ix20084 (.Y (nx20083), .A0 (booth_booth_integration_output_4_9), .A1 (
             nx10266), .S0 (nx36109)) ;
    mux21_ni ix10267 (.Y (nx10266), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_4_10), .S0 (nx36119)) ;
    mux21_ni ix20074 (.Y (nx20073), .A0 (booth_booth_integration_output_4_10), .A1 (
             nx10254), .S0 (nx36111)) ;
    mux21_ni ix10255 (.Y (nx10254), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_4_11), .S0 (nx36119)) ;
    mux21_ni ix20064 (.Y (nx20063), .A0 (booth_booth_integration_output_4_11), .A1 (
             nx10242), .S0 (nx36111)) ;
    mux21_ni ix10243 (.Y (nx10242), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_4_12), .S0 (nx36119)) ;
    mux21_ni ix20054 (.Y (nx20053), .A0 (booth_booth_integration_output_4_12), .A1 (
             nx10230), .S0 (nx36111)) ;
    mux21_ni ix10231 (.Y (nx10230), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_4_13), .S0 (nx36121)) ;
    mux21_ni ix20044 (.Y (nx20043), .A0 (booth_booth_integration_output_4_13), .A1 (
             nx10218), .S0 (nx36111)) ;
    mux21_ni ix10219 (.Y (nx10218), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_4_14), .S0 (nx36121)) ;
    mux21_ni ix20034 (.Y (nx20033), .A0 (booth_booth_integration_output_4_14), .A1 (
             nx10206), .S0 (nx36111)) ;
    mux21_ni ix10207 (.Y (nx10206), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_4_15), .S0 (nx36121)) ;
    mux21 ix20024 (.Y (nx20023), .A0 (nx29480), .A1 (nx29122), .S0 (nx36111)) ;
    mux21_ni ix19674 (.Y (nx19673), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_0), .A1 (nx34939), .S0 (
             nx35823)) ;
    and02 ix19660 (.Y (nx19659), .A0 (nx36349), .A1 (
          booth_booth_integrtaion_4_shift_Reg_count_0)) ;
    mux21_ni ix19854 (.Y (nx19853), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_9), .A1 (nx34925), .S0 (
             nx35823)) ;
    mux21_ni ix19844 (.Y (nx19843), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_8), .S0 (nx36111)) ;
    mux21_ni ix19834 (.Y (nx19833), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_8), .S0 (nx35823)) ;
    mux21_ni ix19824 (.Y (nx19823), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_7), .S0 (nx36113)) ;
    mux21_ni ix19814 (.Y (nx19813), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_7), .S0 (nx35823)) ;
    mux21_ni ix19804 (.Y (nx19803), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_6), .S0 (nx36113)) ;
    mux21_ni ix19794 (.Y (nx19793), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_6), .S0 (nx35823)) ;
    mux21_ni ix19784 (.Y (nx19783), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_5), .S0 (nx36113)) ;
    mux21_ni ix19774 (.Y (nx19773), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_5), .S0 (nx35823)) ;
    mux21_ni ix19764 (.Y (nx19763), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_4), .S0 (nx36113)) ;
    mux21_ni ix19754 (.Y (nx19753), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_4), .S0 (nx35825)) ;
    mux21_ni ix19744 (.Y (nx19743), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_3), .S0 (nx36113)) ;
    mux21_ni ix19734 (.Y (nx19733), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_3), .S0 (nx35825)) ;
    mux21_ni ix19724 (.Y (nx19723), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_2), .S0 (nx36113)) ;
    mux21_ni ix19714 (.Y (nx19713), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_2), .S0 (nx35825)) ;
    mux21_ni ix19704 (.Y (nx19703), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_1), .S0 (nx36113)) ;
    mux21_ni ix19694 (.Y (nx19693), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_4_shift_Reg_output_1), .S0 (nx35825)) ;
    mux21_ni ix19684 (.Y (nx19683), .A0 (
             booth_booth_integrtaion_4_shift_Reg_count_1), .A1 (nx34939), .S0 (
             nx36115)) ;
    and02 ix9647 (.Y (nx9646), .A0 (nx29195), .A1 (nx35763)) ;
    or03 ix29198 (.Y (nx29197), .A0 (nx29199), .A1 (
         booth_booth_integrtaion_4_shift_reg_output_0), .A2 (nx36349)) ;
    mux21_ni ix20014 (.Y (nx20013), .A0 (
             booth_booth_integrtaion_4_booth_output_16), .A1 (nx10176), .S0 (
             nx36115)) ;
    nor02ii ix10177 (.Y (nx10176), .A0 (nx29206), .A1 (nx36121)) ;
    nor02ii ix9653 (.Y (nx9652), .A0 (nx29190), .A1 (
            booth_booth_integrtaion_4_booth_output_16)) ;
    xor2 ix10171 (.Y (nx13217), .A0 (nx29212), .A1 (nx29476)) ;
    xor2 ix10159 (.Y (nx13219), .A0 (nx29237), .A1 (nx35437)) ;
    mux21_ni ix19994 (.Y (nx19993), .A0 (
             booth_booth_integrtaion_4_booth_output_18), .A1 (nx10152), .S0 (
             nx36115)) ;
    nor02ii ix10153 (.Y (nx10152), .A0 (nx29227), .A1 (nx36121)) ;
    xor2 ix10147 (.Y (nx13221), .A0 (nx29242), .A1 (nx29473)) ;
    or02 ix29259 (.Y (nx29258), .A0 (nx29195), .A1 (nx35765)) ;
    xor2 ix10135 (.Y (nx13223), .A0 (nx29276), .A1 (nx35439)) ;
    mux21_ni ix19974 (.Y (nx19973), .A0 (
             booth_booth_integrtaion_4_booth_output_20), .A1 (nx10128), .S0 (
             nx36115)) ;
    nor02ii ix10129 (.Y (nx10128), .A0 (nx29264), .A1 (nx36121)) ;
    xor2 ix10123 (.Y (nx13224), .A0 (nx29281), .A1 (nx29470)) ;
    xor2 ix10111 (.Y (nx13225), .A0 (nx29311), .A1 (nx35441)) ;
    mux21_ni ix19954 (.Y (nx19953), .A0 (
             booth_booth_integrtaion_4_booth_output_22), .A1 (nx10104), .S0 (
             nx36115)) ;
    nor02ii ix10105 (.Y (nx10104), .A0 (nx29299), .A1 (nx36121)) ;
    xor2 ix10099 (.Y (nx13226), .A0 (nx29316), .A1 (nx29467)) ;
    xor2 ix10087 (.Y (nx13227), .A0 (nx29346), .A1 (nx35443)) ;
    mux21_ni ix19934 (.Y (nx19933), .A0 (
             booth_booth_integrtaion_4_booth_output_24), .A1 (nx10080), .S0 (
             nx36115)) ;
    nor02ii ix10081 (.Y (nx10080), .A0 (nx29334), .A1 (nx36123)) ;
    xor2 ix10075 (.Y (nx13228), .A0 (nx29351), .A1 (nx29464)) ;
    xor2 ix10063 (.Y (nx13229), .A0 (nx29381), .A1 (nx35445)) ;
    mux21_ni ix19914 (.Y (nx19913), .A0 (
             booth_booth_integrtaion_4_booth_output_26), .A1 (nx10056), .S0 (
             nx36115)) ;
    nor02ii ix10057 (.Y (nx10056), .A0 (nx29369), .A1 (nx36123)) ;
    xor2 ix10051 (.Y (nx13231), .A0 (nx29386), .A1 (nx29461)) ;
    xor2 ix10039 (.Y (nx13233), .A0 (nx29416), .A1 (nx35447)) ;
    mux21_ni ix19894 (.Y (nx19893), .A0 (
             booth_booth_integrtaion_4_booth_output_28), .A1 (nx10032), .S0 (
             nx35429)) ;
    nor02ii ix10033 (.Y (nx10032), .A0 (nx29404), .A1 (nx36123)) ;
    xor2 ix10027 (.Y (nx13235), .A0 (nx29421), .A1 (nx29458)) ;
    xor2 ix10015 (.Y (nx13236), .A0 (nx29451), .A1 (nx35449)) ;
    mux21_ni ix19874 (.Y (nx19873), .A0 (
             booth_booth_integrtaion_4_booth_output_31), .A1 (nx10008), .S0 (
             nx35429)) ;
    nor02ii ix10009 (.Y (nx10008), .A0 (nx29439), .A1 (nx36123)) ;
    xor2 ix10003 (.Y (nx10002), .A0 (nx29451), .A1 (nx29454)) ;
    nor02ii ix10189 (.Y (nx10188), .A0 (nx9652), .A1 (nx36123)) ;
    and04 ix29499 (.Y (nx29498), .A0 (max_calc_state_0), .A1 (nx35979), .A2 (
          nx35959), .A3 (nx26203)) ;
    mux21_ni ix21034 (.Y (nx21033), .A0 (label_6_output[0]), .A1 (
             label_6_input_0), .S0 (nx36251)) ;
    mux21_ni ix21024 (.Y (nx21023), .A0 (label_6_input_state_machine_0), .A1 (
             mdr_data_out[80]), .S0 (nx36211)) ;
    mux21_ni ix21014 (.Y (nx21013), .A0 (nx35767), .A1 (nx11696), .S0 (nx35479)
             ) ;
    mux21_ni ix11697 (.Y (nx11696), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_5_1), .S0 (nx36139)) ;
    mux21_ni ix21004 (.Y (nx21003), .A0 (booth_booth_integration_output_5_1), .A1 (
             nx11684), .S0 (nx35479)) ;
    mux21_ni ix11685 (.Y (nx11684), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_5_2), .S0 (nx36139)) ;
    mux21_ni ix20994 (.Y (nx20993), .A0 (booth_booth_integration_output_5_2), .A1 (
             nx11672), .S0 (nx35479)) ;
    mux21_ni ix11673 (.Y (nx11672), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_5_3), .S0 (nx36139)) ;
    mux21_ni ix20984 (.Y (nx20983), .A0 (booth_booth_integration_output_5_3), .A1 (
             nx11660), .S0 (nx35479)) ;
    mux21_ni ix11661 (.Y (nx11660), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_5_4), .S0 (nx36139)) ;
    mux21_ni ix20974 (.Y (nx20973), .A0 (booth_booth_integration_output_5_4), .A1 (
             nx11648), .S0 (nx35479)) ;
    mux21_ni ix11649 (.Y (nx11648), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_5_5), .S0 (nx36139)) ;
    mux21_ni ix20964 (.Y (nx20963), .A0 (booth_booth_integration_output_5_5), .A1 (
             nx11636), .S0 (nx35479)) ;
    mux21_ni ix11637 (.Y (nx11636), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_5_6), .S0 (nx36141)) ;
    mux21_ni ix20954 (.Y (nx20953), .A0 (booth_booth_integration_output_5_6), .A1 (
             nx11624), .S0 (nx35479)) ;
    mux21_ni ix11625 (.Y (nx11624), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_5_7), .S0 (nx36141)) ;
    mux21_ni ix20944 (.Y (nx20943), .A0 (booth_booth_integration_output_5_7), .A1 (
             nx11612), .S0 (nx36131)) ;
    mux21_ni ix11613 (.Y (nx11612), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_5_8), .S0 (nx36141)) ;
    mux21_ni ix20934 (.Y (nx20933), .A0 (booth_booth_integration_output_5_8), .A1 (
             nx11600), .S0 (nx36131)) ;
    mux21_ni ix11601 (.Y (nx11600), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_5_9), .S0 (nx36141)) ;
    mux21_ni ix20924 (.Y (nx20923), .A0 (booth_booth_integration_output_5_9), .A1 (
             nx11588), .S0 (nx36131)) ;
    mux21_ni ix11589 (.Y (nx11588), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_5_10), .S0 (nx36141)) ;
    mux21_ni ix20914 (.Y (nx20913), .A0 (booth_booth_integration_output_5_10), .A1 (
             nx11576), .S0 (nx36133)) ;
    mux21_ni ix11577 (.Y (nx11576), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_5_11), .S0 (nx36141)) ;
    mux21_ni ix20904 (.Y (nx20903), .A0 (booth_booth_integration_output_5_11), .A1 (
             nx11564), .S0 (nx36133)) ;
    mux21_ni ix11565 (.Y (nx11564), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_5_12), .S0 (nx36141)) ;
    mux21_ni ix20894 (.Y (nx20893), .A0 (booth_booth_integration_output_5_12), .A1 (
             nx11552), .S0 (nx36133)) ;
    mux21_ni ix11553 (.Y (nx11552), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_5_13), .S0 (nx36143)) ;
    mux21_ni ix20884 (.Y (nx20883), .A0 (booth_booth_integration_output_5_13), .A1 (
             nx11540), .S0 (nx36133)) ;
    mux21_ni ix11541 (.Y (nx11540), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_5_14), .S0 (nx36143)) ;
    mux21_ni ix20874 (.Y (nx20873), .A0 (booth_booth_integration_output_5_14), .A1 (
             nx11528), .S0 (nx36133)) ;
    mux21_ni ix11529 (.Y (nx11528), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_5_15), .S0 (nx36143)) ;
    mux21 ix20864 (.Y (nx20863), .A0 (nx29921), .A1 (nx29563), .S0 (nx36133)) ;
    mux21_ni ix20514 (.Y (nx20513), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_0), .A1 (nx34971), .S0 (
             nx35827)) ;
    and02 ix20500 (.Y (nx20499), .A0 (nx36353), .A1 (
          booth_booth_integrtaion_5_shift_Reg_count_0)) ;
    mux21_ni ix20694 (.Y (nx20693), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_9), .A1 (nx34957), .S0 (
             nx35827)) ;
    mux21_ni ix20684 (.Y (nx20683), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_8), .S0 (nx36133)) ;
    mux21_ni ix20674 (.Y (nx20673), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_8), .S0 (nx35827)) ;
    mux21_ni ix20664 (.Y (nx20663), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_7), .S0 (nx36135)) ;
    mux21_ni ix20654 (.Y (nx20653), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_7), .S0 (nx35827)) ;
    mux21_ni ix20644 (.Y (nx20643), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_6), .S0 (nx36135)) ;
    mux21_ni ix20634 (.Y (nx20633), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_6), .S0 (nx35827)) ;
    mux21_ni ix20624 (.Y (nx20623), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_5), .S0 (nx36135)) ;
    mux21_ni ix20614 (.Y (nx20613), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_5), .S0 (nx35827)) ;
    mux21_ni ix20604 (.Y (nx20603), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_4), .S0 (nx36135)) ;
    mux21_ni ix20594 (.Y (nx20593), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_4), .S0 (nx35829)) ;
    mux21_ni ix20584 (.Y (nx20583), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_3), .S0 (nx36135)) ;
    mux21_ni ix20574 (.Y (nx20573), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_3), .S0 (nx35829)) ;
    mux21_ni ix20564 (.Y (nx20563), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_2), .S0 (nx36135)) ;
    mux21_ni ix20554 (.Y (nx20553), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_2), .S0 (nx35829)) ;
    mux21_ni ix20544 (.Y (nx20543), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_1), .S0 (nx36135)) ;
    mux21_ni ix20534 (.Y (nx20533), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_5_shift_Reg_output_1), .S0 (nx35829)) ;
    mux21_ni ix20524 (.Y (nx20523), .A0 (
             booth_booth_integrtaion_5_shift_Reg_count_1), .A1 (nx34971), .S0 (
             nx36137)) ;
    and02 ix10969 (.Y (nx10968), .A0 (nx29636), .A1 (nx35767)) ;
    or03 ix29639 (.Y (nx29638), .A0 (nx29640), .A1 (
         booth_booth_integrtaion_5_shift_reg_output_0), .A2 (nx36353)) ;
    mux21_ni ix20854 (.Y (nx20853), .A0 (
             booth_booth_integrtaion_5_booth_output_16), .A1 (nx11498), .S0 (
             nx36137)) ;
    nor02ii ix11499 (.Y (nx11498), .A0 (nx29647), .A1 (nx36143)) ;
    nor02ii ix10975 (.Y (nx10974), .A0 (nx29631), .A1 (
            booth_booth_integrtaion_5_booth_output_16)) ;
    xor2 ix11493 (.Y (nx13257), .A0 (nx29653), .A1 (nx29917)) ;
    xor2 ix11481 (.Y (nx13259), .A0 (nx29678), .A1 (nx35485)) ;
    mux21_ni ix20834 (.Y (nx20833), .A0 (
             booth_booth_integrtaion_5_booth_output_18), .A1 (nx11474), .S0 (
             nx36137)) ;
    nor02ii ix11475 (.Y (nx11474), .A0 (nx29668), .A1 (nx36143)) ;
    xor2 ix11469 (.Y (nx13260), .A0 (nx29683), .A1 (nx29914)) ;
    or02 ix29700 (.Y (nx29699), .A0 (nx29636), .A1 (nx35769)) ;
    xor2 ix11457 (.Y (nx13261), .A0 (nx29717), .A1 (nx35487)) ;
    mux21_ni ix20814 (.Y (nx20813), .A0 (
             booth_booth_integrtaion_5_booth_output_20), .A1 (nx11450), .S0 (
             nx36137)) ;
    nor02ii ix11451 (.Y (nx11450), .A0 (nx29705), .A1 (nx36143)) ;
    xor2 ix11445 (.Y (nx13262), .A0 (nx29722), .A1 (nx29911)) ;
    xor2 ix11433 (.Y (nx13263), .A0 (nx29752), .A1 (nx35489)) ;
    mux21_ni ix20794 (.Y (nx20793), .A0 (
             booth_booth_integrtaion_5_booth_output_22), .A1 (nx11426), .S0 (
             nx36137)) ;
    nor02ii ix11427 (.Y (nx11426), .A0 (nx29740), .A1 (nx36143)) ;
    xor2 ix11421 (.Y (nx13264), .A0 (nx29757), .A1 (nx29908)) ;
    xor2 ix11409 (.Y (nx13265), .A0 (nx29787), .A1 (nx35491)) ;
    mux21_ni ix20774 (.Y (nx20773), .A0 (
             booth_booth_integrtaion_5_booth_output_24), .A1 (nx11402), .S0 (
             nx36137)) ;
    nor02ii ix11403 (.Y (nx11402), .A0 (nx29775), .A1 (nx36145)) ;
    xor2 ix11397 (.Y (nx13267), .A0 (nx29792), .A1 (nx29905)) ;
    xor2 ix11385 (.Y (nx13269), .A0 (nx29822), .A1 (nx35493)) ;
    mux21_ni ix20754 (.Y (nx20753), .A0 (
             booth_booth_integrtaion_5_booth_output_26), .A1 (nx11378), .S0 (
             nx36137)) ;
    nor02ii ix11379 (.Y (nx11378), .A0 (nx29810), .A1 (nx36145)) ;
    xor2 ix11373 (.Y (nx13271), .A0 (nx29827), .A1 (nx29902)) ;
    xor2 ix11361 (.Y (nx13272), .A0 (nx29857), .A1 (nx35495)) ;
    mux21_ni ix20734 (.Y (nx20733), .A0 (
             booth_booth_integrtaion_5_booth_output_28), .A1 (nx11354), .S0 (
             nx35477)) ;
    nor02ii ix11355 (.Y (nx11354), .A0 (nx29845), .A1 (nx36145)) ;
    xor2 ix11349 (.Y (nx13273), .A0 (nx29862), .A1 (nx29899)) ;
    xor2 ix11337 (.Y (nx13274), .A0 (nx29892), .A1 (nx35497)) ;
    mux21_ni ix20714 (.Y (nx20713), .A0 (
             booth_booth_integrtaion_5_booth_output_31), .A1 (nx11330), .S0 (
             nx35477)) ;
    nor02ii ix11331 (.Y (nx11330), .A0 (nx29880), .A1 (nx36145)) ;
    xor2 ix11325 (.Y (nx11324), .A0 (nx29892), .A1 (nx29895)) ;
    nor02ii ix11511 (.Y (nx11510), .A0 (nx10974), .A1 (nx36145)) ;
    or03 ix29946 (.Y (nx29945), .A0 (nx30129), .A1 (nx36195), .A2 (nx36069)) ;
    mux21_ni ix21304 (.Y (nx21303), .A0 (label_6_output[14]), .A1 (
             label_6_input_14), .S0 (nx36253)) ;
    mux21_ni ix12155 (.Y (nx12154), .A0 (nx12150), .A1 (
             label_6_input_state_machine_14), .S0 (nx35927)) ;
    mux21_ni ix20484 (.Y (nx20483), .A0 (label_6_input_state_machine_14), .A1 (
             mdr_data_out[94]), .S0 (nx36211)) ;
    mux21_ni ix21294 (.Y (nx21293), .A0 (label_6_output[13]), .A1 (
             label_6_input_13), .S0 (nx36253)) ;
    mux21_ni ix12129 (.Y (nx12128), .A0 (nx12124), .A1 (
             label_6_input_state_machine_13), .S0 (nx35927)) ;
    mux21_ni ix21284 (.Y (nx21283), .A0 (label_6_input_state_machine_13), .A1 (
             mdr_data_out[93]), .S0 (nx36211)) ;
    mux21_ni ix21254 (.Y (nx21253), .A0 (label_6_output[11]), .A1 (
             label_6_input_11), .S0 (nx36251)) ;
    mux21_ni ix12065 (.Y (nx12064), .A0 (nx12060), .A1 (
             label_6_input_state_machine_11), .S0 (nx35927)) ;
    mux21_ni ix21244 (.Y (nx21243), .A0 (label_6_input_state_machine_11), .A1 (
             mdr_data_out[91]), .S0 (nx36211)) ;
    mux21_ni ix21214 (.Y (nx21213), .A0 (label_6_output[9]), .A1 (
             label_6_input_9), .S0 (nx36251)) ;
    mux21_ni ix12001 (.Y (nx12000), .A0 (nx11996), .A1 (
             label_6_input_state_machine_9), .S0 (nx35927)) ;
    mux21_ni ix21204 (.Y (nx21203), .A0 (label_6_input_state_machine_9), .A1 (
             mdr_data_out[89]), .S0 (nx35595)) ;
    mux21_ni ix21174 (.Y (nx21173), .A0 (label_6_output[7]), .A1 (
             label_6_input_7), .S0 (nx36251)) ;
    mux21_ni ix11937 (.Y (nx11936), .A0 (nx11932), .A1 (
             label_6_input_state_machine_7), .S0 (nx35929)) ;
    mux21_ni ix21164 (.Y (nx21163), .A0 (label_6_input_state_machine_7), .A1 (
             mdr_data_out[87]), .S0 (nx36213)) ;
    mux21_ni ix21134 (.Y (nx21133), .A0 (label_6_output[5]), .A1 (
             label_6_input_5), .S0 (nx36251)) ;
    mux21_ni ix11873 (.Y (nx11872), .A0 (nx11868), .A1 (
             label_6_input_state_machine_5), .S0 (nx35929)) ;
    mux21_ni ix21124 (.Y (nx21123), .A0 (label_6_input_state_machine_5), .A1 (
             mdr_data_out[85]), .S0 (nx36213)) ;
    mux21_ni ix21094 (.Y (nx21093), .A0 (label_6_output[3]), .A1 (
             label_6_input_3), .S0 (nx36251)) ;
    mux21_ni ix11809 (.Y (nx11808), .A0 (nx11804), .A1 (
             label_6_input_state_machine_3), .S0 (nx35929)) ;
    mux21_ni ix21084 (.Y (nx21083), .A0 (label_6_input_state_machine_3), .A1 (
             mdr_data_out[83]), .S0 (nx36213)) ;
    mux21_ni ix21054 (.Y (nx21053), .A0 (label_6_output[1]), .A1 (
             label_6_input_1), .S0 (nx36391)) ;
    mux21_ni ix11745 (.Y (nx11744), .A0 (nx11740), .A1 (
             label_6_input_state_machine_1), .S0 (nx35929)) ;
    mux21_ni ix21044 (.Y (nx21043), .A0 (label_6_input_state_machine_1), .A1 (
             mdr_data_out[81]), .S0 (nx36213)) ;
    xnor2 ix30038 (.Y (nx30037), .A0 (nx29935), .A1 (nx30047)) ;
    mux21_ni ix21074 (.Y (nx21073), .A0 (label_6_output[2]), .A1 (
             label_6_input_2), .S0 (nx36391)) ;
    mux21_ni ix11777 (.Y (nx11776), .A0 (nx11772), .A1 (
             label_6_input_state_machine_2), .S0 (nx35929)) ;
    mux21_ni ix21064 (.Y (nx21063), .A0 (label_6_input_state_machine_2), .A1 (
             mdr_data_out[82]), .S0 (nx36213)) ;
    xnor2 ix30053 (.Y (nx30052), .A0 (nx29933), .A1 (nx30062)) ;
    mux21_ni ix21114 (.Y (nx21113), .A0 (label_6_output[4]), .A1 (
             label_6_input_4), .S0 (nx36391)) ;
    mux21_ni ix11841 (.Y (nx11840), .A0 (nx11836), .A1 (
             label_6_input_state_machine_4), .S0 (nx35929)) ;
    mux21_ni ix21104 (.Y (nx21103), .A0 (label_6_input_state_machine_4), .A1 (
             mdr_data_out[84]), .S0 (nx36213)) ;
    xnor2 ix30068 (.Y (nx30067), .A0 (nx29931), .A1 (nx30077)) ;
    mux21_ni ix21154 (.Y (nx21153), .A0 (label_6_output[6]), .A1 (
             label_6_input_6), .S0 (nx36391)) ;
    mux21_ni ix11905 (.Y (nx11904), .A0 (nx11900), .A1 (
             label_6_input_state_machine_6), .S0 (nx35929)) ;
    mux21_ni ix21144 (.Y (nx21143), .A0 (label_6_input_state_machine_6), .A1 (
             mdr_data_out[86]), .S0 (nx36213)) ;
    xnor2 ix30083 (.Y (nx30082), .A0 (nx29929), .A1 (nx30092)) ;
    mux21_ni ix21194 (.Y (nx21193), .A0 (label_6_output[8]), .A1 (
             label_6_input_8), .S0 (nx36391)) ;
    mux21_ni ix11969 (.Y (nx11968), .A0 (nx11964), .A1 (
             label_6_input_state_machine_8), .S0 (nx35931)) ;
    mux21_ni ix21184 (.Y (nx21183), .A0 (label_6_input_state_machine_8), .A1 (
             mdr_data_out[88]), .S0 (nx36215)) ;
    xnor2 ix30098 (.Y (nx30097), .A0 (nx29927), .A1 (nx30107)) ;
    mux21_ni ix21234 (.Y (nx21233), .A0 (label_6_output[10]), .A1 (
             label_6_input_10), .S0 (nx36391)) ;
    mux21_ni ix12033 (.Y (nx12032), .A0 (nx12028), .A1 (
             label_6_input_state_machine_10), .S0 (nx35931)) ;
    mux21_ni ix21224 (.Y (nx21223), .A0 (label_6_input_state_machine_10), .A1 (
             mdr_data_out[90]), .S0 (nx36215)) ;
    xnor2 ix30113 (.Y (nx30112), .A0 (nx29925), .A1 (nx30122)) ;
    mux21_ni ix21274 (.Y (nx21273), .A0 (label_6_output[12]), .A1 (
             label_6_input_12), .S0 (nx36391)) ;
    mux21_ni ix12097 (.Y (nx12096), .A0 (nx12092), .A1 (
             label_6_input_state_machine_12), .S0 (nx35931)) ;
    mux21_ni ix21264 (.Y (nx21263), .A0 (label_6_input_state_machine_12), .A1 (
             mdr_data_out[92]), .S0 (nx36215)) ;
    xnor2 ix30128 (.Y (nx30127), .A0 (nx29923), .A1 (nx30129)) ;
    or03 ix30135 (.Y (nx30134), .A0 (nx30318), .A1 (nx36195), .A2 (nx36069)) ;
    mux21_ni ix20464 (.Y (nx20463), .A0 (label_5_output[14]), .A1 (
             label_5_input_14), .S0 (nx36253)) ;
    mux21_ni ix10833 (.Y (nx10832), .A0 (nx10828), .A1 (
             label_5_input_state_machine_14), .S0 (nx35931)) ;
    mux21_ni ix19644 (.Y (nx19643), .A0 (label_5_input_state_machine_14), .A1 (
             mdr_data_out[78]), .S0 (nx36215)) ;
    mux21_ni ix20454 (.Y (nx20453), .A0 (label_5_output[13]), .A1 (
             label_5_input_13), .S0 (nx36253)) ;
    mux21_ni ix10807 (.Y (nx10806), .A0 (nx10802), .A1 (
             label_5_input_state_machine_13), .S0 (nx35931)) ;
    mux21_ni ix20444 (.Y (nx20443), .A0 (label_5_input_state_machine_13), .A1 (
             mdr_data_out[77]), .S0 (nx36215)) ;
    mux21_ni ix20414 (.Y (nx20413), .A0 (label_5_output[11]), .A1 (
             label_5_input_11), .S0 (nx36253)) ;
    mux21_ni ix10743 (.Y (nx10742), .A0 (nx10738), .A1 (
             label_5_input_state_machine_11), .S0 (nx35931)) ;
    mux21_ni ix20404 (.Y (nx20403), .A0 (label_5_input_state_machine_11), .A1 (
             mdr_data_out[75]), .S0 (nx36215)) ;
    mux21_ni ix20374 (.Y (nx20373), .A0 (label_5_output[9]), .A1 (
             label_5_input_9), .S0 (nx36253)) ;
    mux21_ni ix10679 (.Y (nx10678), .A0 (nx10674), .A1 (
             label_5_input_state_machine_9), .S0 (nx35931)) ;
    mux21_ni ix20364 (.Y (nx20363), .A0 (label_5_input_state_machine_9), .A1 (
             mdr_data_out[73]), .S0 (nx36215)) ;
    mux21_ni ix20334 (.Y (nx20333), .A0 (label_5_output[7]), .A1 (
             label_5_input_7), .S0 (nx36253)) ;
    mux21_ni ix10615 (.Y (nx10614), .A0 (nx10610), .A1 (
             label_5_input_state_machine_7), .S0 (nx35933)) ;
    mux21_ni ix20324 (.Y (nx20323), .A0 (label_5_input_state_machine_7), .A1 (
             mdr_data_out[71]), .S0 (nx36217)) ;
    mux21_ni ix20294 (.Y (nx20293), .A0 (label_5_output[5]), .A1 (
             label_5_input_5), .S0 (nx36255)) ;
    mux21_ni ix10551 (.Y (nx10550), .A0 (nx10546), .A1 (
             label_5_input_state_machine_5), .S0 (nx35933)) ;
    mux21_ni ix20284 (.Y (nx20283), .A0 (label_5_input_state_machine_5), .A1 (
             mdr_data_out[69]), .S0 (nx36217)) ;
    mux21_ni ix20254 (.Y (nx20253), .A0 (label_5_output[3]), .A1 (
             label_5_input_3), .S0 (nx36255)) ;
    mux21_ni ix10487 (.Y (nx10486), .A0 (nx10482), .A1 (
             label_5_input_state_machine_3), .S0 (nx35933)) ;
    mux21_ni ix20244 (.Y (nx20243), .A0 (label_5_input_state_machine_3), .A1 (
             mdr_data_out[67]), .S0 (nx36217)) ;
    mux21_ni ix20214 (.Y (nx20213), .A0 (label_5_output[1]), .A1 (
             label_5_input_1), .S0 (nx36255)) ;
    mux21_ni ix10423 (.Y (nx10422), .A0 (nx10418), .A1 (
             label_5_input_state_machine_1), .S0 (nx35933)) ;
    mux21_ni ix20204 (.Y (nx20203), .A0 (label_5_input_state_machine_1), .A1 (
             mdr_data_out[65]), .S0 (nx36217)) ;
    xnor2 ix30227 (.Y (nx30226), .A0 (nx29494), .A1 (nx30236)) ;
    mux21_ni ix20234 (.Y (nx20233), .A0 (label_5_output[2]), .A1 (
             label_5_input_2), .S0 (nx36255)) ;
    mux21_ni ix10455 (.Y (nx10454), .A0 (nx10450), .A1 (
             label_5_input_state_machine_2), .S0 (nx35933)) ;
    mux21_ni ix20224 (.Y (nx20223), .A0 (label_5_input_state_machine_2), .A1 (
             mdr_data_out[66]), .S0 (nx36217)) ;
    xnor2 ix30242 (.Y (nx30241), .A0 (nx29492), .A1 (nx30251)) ;
    mux21_ni ix20274 (.Y (nx20273), .A0 (label_5_output[4]), .A1 (
             label_5_input_4), .S0 (nx36255)) ;
    mux21_ni ix10519 (.Y (nx10518), .A0 (nx10514), .A1 (
             label_5_input_state_machine_4), .S0 (nx35933)) ;
    mux21_ni ix20264 (.Y (nx20263), .A0 (label_5_input_state_machine_4), .A1 (
             mdr_data_out[68]), .S0 (nx36217)) ;
    xnor2 ix30257 (.Y (nx30256), .A0 (nx29490), .A1 (nx30266)) ;
    mux21_ni ix20314 (.Y (nx20313), .A0 (label_5_output[6]), .A1 (
             label_5_input_6), .S0 (nx36255)) ;
    mux21_ni ix10583 (.Y (nx10582), .A0 (nx10578), .A1 (
             label_5_input_state_machine_6), .S0 (nx35933)) ;
    mux21_ni ix20304 (.Y (nx20303), .A0 (label_5_input_state_machine_6), .A1 (
             mdr_data_out[70]), .S0 (nx36217)) ;
    xnor2 ix30272 (.Y (nx30271), .A0 (nx29488), .A1 (nx30281)) ;
    mux21_ni ix20354 (.Y (nx20353), .A0 (label_5_output[8]), .A1 (
             label_5_input_8), .S0 (nx36255)) ;
    mux21_ni ix10647 (.Y (nx10646), .A0 (nx10642), .A1 (
             label_5_input_state_machine_8), .S0 (nx35935)) ;
    mux21_ni ix20344 (.Y (nx20343), .A0 (label_5_input_state_machine_8), .A1 (
             mdr_data_out[72]), .S0 (nx36219)) ;
    xnor2 ix30287 (.Y (nx30286), .A0 (nx29486), .A1 (nx30296)) ;
    mux21_ni ix20394 (.Y (nx20393), .A0 (label_5_output[10]), .A1 (
             label_5_input_10), .S0 (nx36257)) ;
    mux21_ni ix10711 (.Y (nx10710), .A0 (nx10706), .A1 (
             label_5_input_state_machine_10), .S0 (nx35935)) ;
    mux21_ni ix20384 (.Y (nx20383), .A0 (label_5_input_state_machine_10), .A1 (
             mdr_data_out[74]), .S0 (nx36219)) ;
    xnor2 ix30302 (.Y (nx30301), .A0 (nx29484), .A1 (nx30311)) ;
    mux21_ni ix20434 (.Y (nx20433), .A0 (label_5_output[12]), .A1 (
             label_5_input_12), .S0 (nx36257)) ;
    mux21_ni ix10775 (.Y (nx10774), .A0 (nx10770), .A1 (
             label_5_input_state_machine_12), .S0 (nx35935)) ;
    mux21_ni ix20424 (.Y (nx20423), .A0 (label_5_input_state_machine_12), .A1 (
             mdr_data_out[76]), .S0 (nx36219)) ;
    xnor2 ix30317 (.Y (nx30316), .A0 (nx29482), .A1 (nx30318)) ;
    xnor2 ix12177 (.Y (nx12176), .A0 (nx29942), .A1 (nx30132)) ;
    xnor2 ix30322 (.Y (nx30321), .A0 (nx30325), .A1 (
          max_calc_comparator_third_inp1_13)) ;
    or03 ix30340 (.Y (nx30339), .A0 (nx30122), .A1 (nx36197), .A2 (nx36069)) ;
    or03 ix30346 (.Y (nx30345), .A0 (nx30311), .A1 (nx36197), .A2 (nx36069)) ;
    xnor2 ix12221 (.Y (nx12220), .A0 (nx30336), .A1 (nx30343)) ;
    xnor2 ix30350 (.Y (nx30349), .A0 (nx30353), .A1 (
          max_calc_comparator_third_inp1_11)) ;
    or03 ix30368 (.Y (nx30367), .A0 (nx30107), .A1 (nx36197), .A2 (nx36069)) ;
    or03 ix30374 (.Y (nx30373), .A0 (nx30296), .A1 (nx36197), .A2 (nx36069)) ;
    xnor2 ix12265 (.Y (nx12264), .A0 (nx30364), .A1 (nx30371)) ;
    xnor2 ix30378 (.Y (nx30377), .A0 (nx30381), .A1 (
          max_calc_comparator_third_inp1_9)) ;
    or03 ix30396 (.Y (nx30395), .A0 (nx30092), .A1 (nx36197), .A2 (nx36069)) ;
    or03 ix30402 (.Y (nx30401), .A0 (nx30281), .A1 (nx36197), .A2 (nx35365)) ;
    xnor2 ix12309 (.Y (nx12308), .A0 (nx30392), .A1 (nx30399)) ;
    xnor2 ix30406 (.Y (nx30405), .A0 (nx30409), .A1 (
          max_calc_comparator_third_inp1_7)) ;
    or03 ix30424 (.Y (nx30423), .A0 (nx30077), .A1 (nx36197), .A2 (nx35365)) ;
    or03 ix30430 (.Y (nx30429), .A0 (nx30266), .A1 (nx36199), .A2 (nx35365)) ;
    xnor2 ix12353 (.Y (nx12352), .A0 (nx30420), .A1 (nx30427)) ;
    xnor2 ix30434 (.Y (nx30433), .A0 (nx30437), .A1 (
          max_calc_comparator_third_inp1_5)) ;
    or03 ix30452 (.Y (nx30451), .A0 (nx30062), .A1 (nx36199), .A2 (nx35365)) ;
    or03 ix30458 (.Y (nx30457), .A0 (nx30251), .A1 (nx36199), .A2 (nx35365)) ;
    xnor2 ix12397 (.Y (nx12396), .A0 (nx30448), .A1 (nx30455)) ;
    xnor2 ix30462 (.Y (nx30461), .A0 (nx30465), .A1 (
          max_calc_comparator_third_inp1_3)) ;
    or03 ix30480 (.Y (nx30479), .A0 (nx30047), .A1 (nx36199), .A2 (nx35365)) ;
    or03 ix30486 (.Y (nx30485), .A0 (nx30236), .A1 (nx36199), .A2 (nx36073)) ;
    xnor2 ix12441 (.Y (nx12440), .A0 (nx30476), .A1 (nx30483)) ;
    xnor2 ix12463 (.Y (nx12462), .A0 (nx30491), .A1 (nx30495)) ;
    xnor2 ix12689 (.Y (nx12688), .A0 (nx30506), .A1 (nx30524)) ;
    mux21_ni ix21614 (.Y (nx21613), .A0 (label_6_output[15]), .A1 (
             label_6_input_15), .S0 (nx36257)) ;
    mux21_ni ix12625 (.Y (nx12624), .A0 (nx12620), .A1 (
             label_6_input_state_machine_15), .S0 (nx35935)) ;
    mux21_ni ix21604 (.Y (nx21603), .A0 (label_6_input_state_machine_15), .A1 (
             mdr_data_out[95]), .S0 (nx36219)) ;
    xor2 ix30520 (.Y (nx30519), .A0 (nx29921), .A1 (label_6_output[15])) ;
    mux21_ni ix21644 (.Y (nx21643), .A0 (label_5_output[15]), .A1 (
             label_5_input_15), .S0 (nx36257)) ;
    mux21_ni ix12667 (.Y (nx12666), .A0 (nx12662), .A1 (
             label_5_input_state_machine_15), .S0 (nx35935)) ;
    mux21_ni ix21634 (.Y (nx21633), .A0 (label_5_input_state_machine_15), .A1 (
             mdr_data_out[79]), .S0 (nx36219)) ;
    xor2 ix30538 (.Y (nx30537), .A0 (nx29480), .A1 (label_5_output[15])) ;
    nand02 ix9537 (.Y (nx34913), .A0 (nx36291), .A1 (nx35869)) ;
    nand04 ix9533 (.Y (nx34905), .A0 (nx36291), .A1 (nx35737), .A2 (nx26203), .A3 (
           nx35641)) ;
    mux21_ni ix16897 (.Y (nx16896), .A0 (max_calc_ans4_0), .A1 (
             label_4_output[0]), .S0 (nx35979)) ;
    mux21_ni ix14674 (.Y (nx14673), .A0 (label_4_output[0]), .A1 (
             label_4_input_0), .S0 (nx36257)) ;
    mux21_ni ix14664 (.Y (nx14663), .A0 (label_4_input_state_machine_0), .A1 (
             mdr_data_out[48]), .S0 (nx36219)) ;
    mux21_ni ix14654 (.Y (nx14653), .A0 (nx35719), .A1 (nx1722), .S0 (nx35505)
             ) ;
    mux21_ni ix1723 (.Y (nx1722), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_3_1), .S0 (nx36155)) ;
    mux21_ni ix14644 (.Y (nx14643), .A0 (booth_booth_integration_output_3_1), .A1 (
             nx1710), .S0 (nx35505)) ;
    mux21_ni ix1711 (.Y (nx1710), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_3_2), .S0 (nx36155)) ;
    mux21_ni ix14634 (.Y (nx14633), .A0 (booth_booth_integration_output_3_2), .A1 (
             nx1698), .S0 (nx35505)) ;
    mux21_ni ix1699 (.Y (nx1698), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_3_3), .S0 (nx36155)) ;
    mux21_ni ix14624 (.Y (nx14623), .A0 (booth_booth_integration_output_3_3), .A1 (
             nx1686), .S0 (nx35505)) ;
    mux21_ni ix1687 (.Y (nx1686), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_3_4), .S0 (nx36155)) ;
    mux21_ni ix14614 (.Y (nx14613), .A0 (booth_booth_integration_output_3_4), .A1 (
             nx1674), .S0 (nx35505)) ;
    mux21_ni ix1675 (.Y (nx1674), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_3_5), .S0 (nx36155)) ;
    mux21_ni ix14604 (.Y (nx14603), .A0 (booth_booth_integration_output_3_5), .A1 (
             nx1662), .S0 (nx35505)) ;
    mux21_ni ix1663 (.Y (nx1662), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_3_6), .S0 (nx36157)) ;
    mux21_ni ix14594 (.Y (nx14593), .A0 (booth_booth_integration_output_3_6), .A1 (
             nx1650), .S0 (nx35505)) ;
    mux21_ni ix1651 (.Y (nx1650), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_3_7), .S0 (nx36157)) ;
    mux21_ni ix14584 (.Y (nx14583), .A0 (booth_booth_integration_output_3_7), .A1 (
             nx1638), .S0 (nx36147)) ;
    mux21_ni ix1639 (.Y (nx1638), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_3_8), .S0 (nx36157)) ;
    mux21_ni ix14574 (.Y (nx14573), .A0 (booth_booth_integration_output_3_8), .A1 (
             nx1626), .S0 (nx36147)) ;
    mux21_ni ix1627 (.Y (nx1626), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_3_9), .S0 (nx36157)) ;
    mux21_ni ix14564 (.Y (nx14563), .A0 (booth_booth_integration_output_3_9), .A1 (
             nx1614), .S0 (nx36147)) ;
    mux21_ni ix1615 (.Y (nx1614), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_3_10), .S0 (nx36157)) ;
    mux21_ni ix14554 (.Y (nx14553), .A0 (booth_booth_integration_output_3_10), .A1 (
             nx1602), .S0 (nx36149)) ;
    mux21_ni ix1603 (.Y (nx1602), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_3_11), .S0 (nx36157)) ;
    mux21_ni ix14544 (.Y (nx14543), .A0 (booth_booth_integration_output_3_11), .A1 (
             nx1590), .S0 (nx36149)) ;
    mux21_ni ix1591 (.Y (nx1590), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_3_12), .S0 (nx36157)) ;
    mux21_ni ix14534 (.Y (nx14533), .A0 (booth_booth_integration_output_3_12), .A1 (
             nx1578), .S0 (nx36149)) ;
    mux21_ni ix1579 (.Y (nx1578), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_3_13), .S0 (nx36159)) ;
    mux21_ni ix14524 (.Y (nx14523), .A0 (booth_booth_integration_output_3_13), .A1 (
             nx1566), .S0 (nx36149)) ;
    mux21_ni ix1567 (.Y (nx1566), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_3_14), .S0 (nx36159)) ;
    mux21_ni ix14514 (.Y (nx14513), .A0 (booth_booth_integration_output_3_14), .A1 (
             nx1554), .S0 (nx36149)) ;
    mux21_ni ix1555 (.Y (nx1554), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_3_15), .S0 (nx36159)) ;
    mux21 ix14504 (.Y (nx14503), .A0 (nx30966), .A1 (nx30608), .S0 (nx36149)) ;
    mux21_ni ix14154 (.Y (nx14153), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_0), .A1 (nx34571), .S0 (
             nx35831)) ;
    and02 ix14140 (.Y (nx14139), .A0 (nx36315), .A1 (
          booth_booth_integrtaion_3_shift_Reg_count_0)) ;
    mux21_ni ix14334 (.Y (nx14333), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_9), .A1 (nx34557), .S0 (
             nx35831)) ;
    mux21_ni ix14324 (.Y (nx14323), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_8), .S0 (nx36149)) ;
    mux21_ni ix14314 (.Y (nx14313), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_8), .S0 (nx35831)) ;
    mux21_ni ix14304 (.Y (nx14303), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_7), .S0 (nx36151)) ;
    mux21_ni ix14294 (.Y (nx14293), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_7), .S0 (nx35831)) ;
    mux21_ni ix14284 (.Y (nx14283), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_6), .S0 (nx36151)) ;
    mux21_ni ix14274 (.Y (nx14273), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_6), .S0 (nx35831)) ;
    mux21_ni ix14264 (.Y (nx14263), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_5), .S0 (nx36151)) ;
    mux21_ni ix14254 (.Y (nx14253), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_5), .S0 (nx35831)) ;
    mux21_ni ix14244 (.Y (nx14243), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_4), .S0 (nx36151)) ;
    mux21_ni ix14234 (.Y (nx14233), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_4), .S0 (nx35833)) ;
    mux21_ni ix14224 (.Y (nx14223), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_3), .S0 (nx36151)) ;
    mux21_ni ix14214 (.Y (nx14213), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_3), .S0 (nx35833)) ;
    mux21_ni ix14204 (.Y (nx14203), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_2), .S0 (nx36151)) ;
    mux21_ni ix14194 (.Y (nx14193), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_2), .S0 (nx35833)) ;
    mux21_ni ix14184 (.Y (nx14183), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_1), .S0 (nx36151)) ;
    mux21_ni ix14174 (.Y (nx14173), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_3_shift_Reg_output_1), .S0 (nx35833)) ;
    mux21_ni ix14164 (.Y (nx14163), .A0 (
             booth_booth_integrtaion_3_shift_Reg_count_1), .A1 (nx34571), .S0 (
             nx36153)) ;
    and02 ix995 (.Y (nx994), .A0 (nx30681), .A1 (nx35719)) ;
    or03 ix30684 (.Y (nx30683), .A0 (nx30685), .A1 (
         booth_booth_integrtaion_3_shift_reg_output_0), .A2 (nx36315)) ;
    mux21_ni ix14494 (.Y (nx14493), .A0 (
             booth_booth_integrtaion_3_booth_output_16), .A1 (nx1524), .S0 (
             nx36153)) ;
    nor02ii ix1525 (.Y (nx1524), .A0 (nx30692), .A1 (nx36159)) ;
    nor02ii ix1001 (.Y (nx1000), .A0 (nx30676), .A1 (
            booth_booth_integrtaion_3_booth_output_16)) ;
    xor2 ix1519 (.Y (nx12913), .A0 (nx30698), .A1 (nx30962)) ;
    xor2 ix1507 (.Y (nx12915), .A0 (nx30723), .A1 (nx35511)) ;
    mux21_ni ix14474 (.Y (nx14473), .A0 (
             booth_booth_integrtaion_3_booth_output_18), .A1 (nx1500), .S0 (
             nx36153)) ;
    nor02ii ix1501 (.Y (nx1500), .A0 (nx30713), .A1 (nx36159)) ;
    xor2 ix1495 (.Y (nx12917), .A0 (nx30728), .A1 (nx30959)) ;
    or02 ix30745 (.Y (nx30744), .A0 (nx30681), .A1 (nx35721)) ;
    xor2 ix1483 (.Y (nx12919), .A0 (nx30762), .A1 (nx35513)) ;
    mux21_ni ix14454 (.Y (nx14453), .A0 (
             booth_booth_integrtaion_3_booth_output_20), .A1 (nx1476), .S0 (
             nx36153)) ;
    nor02ii ix1477 (.Y (nx1476), .A0 (nx30750), .A1 (nx36159)) ;
    xor2 ix1471 (.Y (nx12921), .A0 (nx30767), .A1 (nx30956)) ;
    xor2 ix1459 (.Y (nx12922), .A0 (nx30797), .A1 (nx35515)) ;
    mux21_ni ix14434 (.Y (nx14433), .A0 (
             booth_booth_integrtaion_3_booth_output_22), .A1 (nx1452), .S0 (
             nx36153)) ;
    nor02ii ix1453 (.Y (nx1452), .A0 (nx30785), .A1 (nx36159)) ;
    xor2 ix1447 (.Y (nx12923), .A0 (nx30802), .A1 (nx30953)) ;
    xor2 ix1435 (.Y (nx12925), .A0 (nx30832), .A1 (nx35517)) ;
    mux21_ni ix14414 (.Y (nx14413), .A0 (
             booth_booth_integrtaion_3_booth_output_24), .A1 (nx1428), .S0 (
             nx36153)) ;
    nor02ii ix1429 (.Y (nx1428), .A0 (nx30820), .A1 (nx36161)) ;
    xor2 ix1423 (.Y (nx12927), .A0 (nx30837), .A1 (nx30950)) ;
    xor2 ix1411 (.Y (nx12929), .A0 (nx30867), .A1 (nx35519)) ;
    mux21_ni ix14394 (.Y (nx14393), .A0 (
             booth_booth_integrtaion_3_booth_output_26), .A1 (nx1404), .S0 (
             nx36153)) ;
    nor02ii ix1405 (.Y (nx1404), .A0 (nx30855), .A1 (nx36161)) ;
    xor2 ix1399 (.Y (nx12930), .A0 (nx30872), .A1 (nx30947)) ;
    xor2 ix1387 (.Y (nx12931), .A0 (nx30902), .A1 (nx35521)) ;
    mux21_ni ix14374 (.Y (nx14373), .A0 (
             booth_booth_integrtaion_3_booth_output_28), .A1 (nx1380), .S0 (
             nx35503)) ;
    nor02ii ix1381 (.Y (nx1380), .A0 (nx30890), .A1 (nx36161)) ;
    xor2 ix1375 (.Y (nx12933), .A0 (nx30907), .A1 (nx30944)) ;
    xor2 ix1363 (.Y (nx12935), .A0 (nx30937), .A1 (nx35523)) ;
    mux21_ni ix14354 (.Y (nx14353), .A0 (
             booth_booth_integrtaion_3_booth_output_31), .A1 (nx1356), .S0 (
             nx35503)) ;
    nor02ii ix1357 (.Y (nx1356), .A0 (nx30925), .A1 (nx36161)) ;
    xor2 ix1351 (.Y (nx1350), .A0 (nx30937), .A1 (nx30940)) ;
    nor02ii ix1537 (.Y (nx1536), .A0 (nx1000), .A1 (nx36161)) ;
    ao32 ix24244 (.Y (nx24243), .A0 (nx35961), .A1 (nx35647), .A2 (nx36291), .B0 (
         max_calc_ans4_0), .B1 (nx35877)) ;
    mux21 ix30987 (.Y (nx35647), .A0 (nx31429), .A1 (nx30990), .S0 (nx35893)) ;
    mux21_ni ix22234 (.Y (nx22233), .A0 (label_7_output[0]), .A1 (
             label_7_input_0), .S0 (nx36257)) ;
    mux21_ni ix22224 (.Y (nx22223), .A0 (label_7_input_state_machine_0), .A1 (
             mdr_data_out[96]), .S0 (nx36219)) ;
    mux21_ni ix22214 (.Y (nx22213), .A0 (nx35771), .A1 (nx13564), .S0 (nx35531)
             ) ;
    mux21_ni ix13565 (.Y (nx13564), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_6_1), .S0 (nx36171)) ;
    mux21_ni ix22204 (.Y (nx22203), .A0 (booth_booth_integration_output_6_1), .A1 (
             nx13552), .S0 (nx35531)) ;
    mux21_ni ix13553 (.Y (nx13552), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_6_2), .S0 (nx36171)) ;
    mux21_ni ix22194 (.Y (nx22193), .A0 (booth_booth_integration_output_6_2), .A1 (
             nx13540), .S0 (nx35531)) ;
    mux21_ni ix13541 (.Y (nx13540), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_6_3), .S0 (nx36171)) ;
    mux21_ni ix22184 (.Y (nx22183), .A0 (booth_booth_integration_output_6_3), .A1 (
             nx13528), .S0 (nx35531)) ;
    mux21_ni ix13529 (.Y (nx13528), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_6_4), .S0 (nx36171)) ;
    mux21_ni ix22174 (.Y (nx22173), .A0 (booth_booth_integration_output_6_4), .A1 (
             nx13516), .S0 (nx35531)) ;
    mux21_ni ix13517 (.Y (nx13516), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_6_5), .S0 (nx36171)) ;
    mux21_ni ix22164 (.Y (nx22163), .A0 (booth_booth_integration_output_6_5), .A1 (
             nx13504), .S0 (nx35531)) ;
    mux21_ni ix13505 (.Y (nx13504), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_6_6), .S0 (nx36173)) ;
    mux21_ni ix22154 (.Y (nx22153), .A0 (booth_booth_integration_output_6_6), .A1 (
             nx13492), .S0 (nx35531)) ;
    mux21_ni ix13493 (.Y (nx13492), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_6_7), .S0 (nx36173)) ;
    mux21_ni ix22144 (.Y (nx22143), .A0 (booth_booth_integration_output_6_7), .A1 (
             nx13480), .S0 (nx36163)) ;
    mux21_ni ix13481 (.Y (nx13480), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_6_8), .S0 (nx36173)) ;
    mux21_ni ix22134 (.Y (nx22133), .A0 (booth_booth_integration_output_6_8), .A1 (
             nx13468), .S0 (nx36163)) ;
    mux21_ni ix13469 (.Y (nx13468), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_6_9), .S0 (nx36173)) ;
    mux21_ni ix22124 (.Y (nx22123), .A0 (booth_booth_integration_output_6_9), .A1 (
             nx13456), .S0 (nx36163)) ;
    mux21_ni ix13457 (.Y (nx13456), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_6_10), .S0 (nx36173)) ;
    mux21_ni ix22114 (.Y (nx22113), .A0 (booth_booth_integration_output_6_10), .A1 (
             nx13444), .S0 (nx36165)) ;
    mux21_ni ix13445 (.Y (nx13444), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_6_11), .S0 (nx36173)) ;
    mux21_ni ix22104 (.Y (nx22103), .A0 (booth_booth_integration_output_6_11), .A1 (
             nx13432), .S0 (nx36165)) ;
    mux21_ni ix13433 (.Y (nx13432), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_6_12), .S0 (nx36173)) ;
    mux21_ni ix22094 (.Y (nx22093), .A0 (booth_booth_integration_output_6_12), .A1 (
             nx13420), .S0 (nx36165)) ;
    mux21_ni ix13421 (.Y (nx13420), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_6_13), .S0 (nx36175)) ;
    mux21_ni ix22084 (.Y (nx22083), .A0 (booth_booth_integration_output_6_13), .A1 (
             nx13408), .S0 (nx36165)) ;
    mux21_ni ix13409 (.Y (nx13408), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_6_14), .S0 (nx36175)) ;
    mux21_ni ix22074 (.Y (nx22073), .A0 (booth_booth_integration_output_6_14), .A1 (
             nx13396), .S0 (nx36165)) ;
    mux21_ni ix13397 (.Y (nx13396), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_6_15), .S0 (nx36175)) ;
    mux21 ix22064 (.Y (nx22063), .A0 (nx31409), .A1 (nx31051), .S0 (nx36165)) ;
    mux21_ni ix21714 (.Y (nx21713), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_0), .A1 (nx35011), .S0 (
             nx35835)) ;
    and02 ix21700 (.Y (nx21699), .A0 (nx36357), .A1 (
          booth_booth_integrtaion_6_shift_Reg_count_0)) ;
    mux21_ni ix21894 (.Y (nx21893), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_9), .A1 (nx34997), .S0 (
             nx35835)) ;
    mux21_ni ix21884 (.Y (nx21883), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_8), .S0 (nx36165)) ;
    mux21_ni ix21874 (.Y (nx21873), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_8), .S0 (nx35835)) ;
    mux21_ni ix21864 (.Y (nx21863), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_7), .S0 (nx36167)) ;
    mux21_ni ix21854 (.Y (nx21853), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_7), .S0 (nx35835)) ;
    mux21_ni ix21844 (.Y (nx21843), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_6), .S0 (nx36167)) ;
    mux21_ni ix21834 (.Y (nx21833), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_6), .S0 (nx35835)) ;
    mux21_ni ix21824 (.Y (nx21823), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_5), .S0 (nx36167)) ;
    mux21_ni ix21814 (.Y (nx21813), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_5), .S0 (nx35835)) ;
    mux21_ni ix21804 (.Y (nx21803), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_4), .S0 (nx36167)) ;
    mux21_ni ix21794 (.Y (nx21793), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_4), .S0 (nx35837)) ;
    mux21_ni ix21784 (.Y (nx21783), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_3), .S0 (nx36167)) ;
    mux21_ni ix21774 (.Y (nx21773), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_3), .S0 (nx35837)) ;
    mux21_ni ix21764 (.Y (nx21763), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_2), .S0 (nx36167)) ;
    mux21_ni ix21754 (.Y (nx21753), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_2), .S0 (nx35837)) ;
    mux21_ni ix21744 (.Y (nx21743), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_1), .S0 (nx36167)) ;
    mux21_ni ix21734 (.Y (nx21733), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_6_shift_Reg_output_1), .S0 (nx35837)) ;
    mux21_ni ix21724 (.Y (nx21723), .A0 (
             booth_booth_integrtaion_6_shift_Reg_count_1), .A1 (nx35011), .S0 (
             nx36169)) ;
    and02 ix12837 (.Y (nx12836), .A0 (nx31124), .A1 (nx35771)) ;
    or03 ix31127 (.Y (nx31126), .A0 (nx31128), .A1 (
         booth_booth_integrtaion_6_shift_reg_output_0), .A2 (nx36357)) ;
    mux21_ni ix22054 (.Y (nx22053), .A0 (
             booth_booth_integrtaion_6_booth_output_16), .A1 (nx13366), .S0 (
             nx36169)) ;
    nor02ii ix13367 (.Y (nx13366), .A0 (nx31135), .A1 (nx36175)) ;
    nor02ii ix12843 (.Y (nx12842), .A0 (nx31119), .A1 (
            booth_booth_integrtaion_6_booth_output_16)) ;
    xor2 ix13361 (.Y (nx13296), .A0 (nx31141), .A1 (nx31405)) ;
    xor2 ix13349 (.Y (nx13297), .A0 (nx31166), .A1 (nx35537)) ;
    mux21_ni ix22034 (.Y (nx22033), .A0 (
             booth_booth_integrtaion_6_booth_output_18), .A1 (nx13342), .S0 (
             nx36169)) ;
    nor02ii ix13343 (.Y (nx13342), .A0 (nx31156), .A1 (nx36175)) ;
    xor2 ix13337 (.Y (nx13298), .A0 (nx31171), .A1 (nx31402)) ;
    or02 ix31188 (.Y (nx31187), .A0 (nx31124), .A1 (nx35773)) ;
    xor2 ix13325 (.Y (nx13299), .A0 (nx31205), .A1 (nx35539)) ;
    mux21_ni ix22014 (.Y (nx22013), .A0 (
             booth_booth_integrtaion_6_booth_output_20), .A1 (nx13318), .S0 (
             nx36169)) ;
    nor02ii ix13319 (.Y (nx13318), .A0 (nx31193), .A1 (nx36175)) ;
    xor2 ix13313 (.Y (nx13300), .A0 (nx31210), .A1 (nx31399)) ;
    xor2 ix13301 (.Y (nx13301), .A0 (nx31240), .A1 (nx35541)) ;
    mux21_ni ix21994 (.Y (nx21993), .A0 (
             booth_booth_integrtaion_6_booth_output_22), .A1 (nx13294), .S0 (
             nx36169)) ;
    nor02ii ix13295 (.Y (nx13294), .A0 (nx31228), .A1 (nx36175)) ;
    xor2 ix13289 (.Y (nx13303), .A0 (nx31245), .A1 (nx31396)) ;
    xor2 ix13277 (.Y (nx13305), .A0 (nx31275), .A1 (nx35543)) ;
    mux21_ni ix21974 (.Y (nx21973), .A0 (
             booth_booth_integrtaion_6_booth_output_24), .A1 (nx13270), .S0 (
             nx36169)) ;
    nor02ii ix13271 (.Y (nx13270), .A0 (nx31263), .A1 (nx36177)) ;
    xor2 ix13265 (.Y (nx13307), .A0 (nx31280), .A1 (nx31393)) ;
    xor2 ix13253 (.Y (nx13308), .A0 (nx31310), .A1 (nx35545)) ;
    mux21_ni ix21954 (.Y (nx21953), .A0 (
             booth_booth_integrtaion_6_booth_output_26), .A1 (nx13246), .S0 (
             nx36169)) ;
    nor02ii ix13247 (.Y (nx13246), .A0 (nx31298), .A1 (nx36177)) ;
    xor2 ix13241 (.Y (nx13309), .A0 (nx31315), .A1 (nx31390)) ;
    xor2 ix13229 (.Y (nx13310), .A0 (nx31345), .A1 (nx35547)) ;
    mux21_ni ix21934 (.Y (nx21933), .A0 (
             booth_booth_integrtaion_6_booth_output_28), .A1 (nx13222), .S0 (
             nx35529)) ;
    nor02ii ix13223 (.Y (nx13222), .A0 (nx31333), .A1 (nx36177)) ;
    xor2 ix13217 (.Y (nx13311), .A0 (nx31350), .A1 (nx31387)) ;
    xor2 ix13205 (.Y (nx13312), .A0 (nx31380), .A1 (nx35549)) ;
    mux21_ni ix21914 (.Y (nx21913), .A0 (
             booth_booth_integrtaion_6_booth_output_31), .A1 (nx13198), .S0 (
             nx35529)) ;
    nor02ii ix13199 (.Y (nx13198), .A0 (nx31368), .A1 (nx36177)) ;
    xor2 ix13193 (.Y (nx13192), .A0 (nx31380), .A1 (nx31383)) ;
    nor02ii ix13379 (.Y (nx13378), .A0 (nx12842), .A1 (nx36177)) ;
    mux21_ni ix23074 (.Y (nx23073), .A0 (label_8_output[0]), .A1 (
             label_8_input_0), .S0 (nx36257)) ;
    mux21_ni ix23064 (.Y (nx23063), .A0 (label_8_input_state_machine_0), .A1 (
             mdr_data_out[112]), .S0 (nx36221)) ;
    mux21_ni ix23054 (.Y (nx23053), .A0 (nx35775), .A1 (nx14880), .S0 (nx35557)
             ) ;
    mux21_ni ix14881 (.Y (nx14880), .A0 (mdr_data_out[0]), .A1 (
             booth_booth_integration_output_7_1), .S0 (nx36187)) ;
    mux21_ni ix23044 (.Y (nx23043), .A0 (booth_booth_integration_output_7_1), .A1 (
             nx14868), .S0 (nx35557)) ;
    mux21_ni ix14869 (.Y (nx14868), .A0 (mdr_data_out[1]), .A1 (
             booth_booth_integration_output_7_2), .S0 (nx36187)) ;
    mux21_ni ix23034 (.Y (nx23033), .A0 (booth_booth_integration_output_7_2), .A1 (
             nx14856), .S0 (nx35557)) ;
    mux21_ni ix14857 (.Y (nx14856), .A0 (mdr_data_out[2]), .A1 (
             booth_booth_integration_output_7_3), .S0 (nx36187)) ;
    mux21_ni ix23024 (.Y (nx23023), .A0 (booth_booth_integration_output_7_3), .A1 (
             nx14844), .S0 (nx35557)) ;
    mux21_ni ix14845 (.Y (nx14844), .A0 (mdr_data_out[3]), .A1 (
             booth_booth_integration_output_7_4), .S0 (nx36187)) ;
    mux21_ni ix23014 (.Y (nx23013), .A0 (booth_booth_integration_output_7_4), .A1 (
             nx14832), .S0 (nx35557)) ;
    mux21_ni ix14833 (.Y (nx14832), .A0 (mdr_data_out[4]), .A1 (
             booth_booth_integration_output_7_5), .S0 (nx36187)) ;
    mux21_ni ix23004 (.Y (nx23003), .A0 (booth_booth_integration_output_7_5), .A1 (
             nx14820), .S0 (nx35557)) ;
    mux21_ni ix14821 (.Y (nx14820), .A0 (mdr_data_out[5]), .A1 (
             booth_booth_integration_output_7_6), .S0 (nx36189)) ;
    mux21_ni ix22994 (.Y (nx22993), .A0 (booth_booth_integration_output_7_6), .A1 (
             nx14808), .S0 (nx35557)) ;
    mux21_ni ix14809 (.Y (nx14808), .A0 (mdr_data_out[6]), .A1 (
             booth_booth_integration_output_7_7), .S0 (nx36189)) ;
    mux21_ni ix22984 (.Y (nx22983), .A0 (booth_booth_integration_output_7_7), .A1 (
             nx14796), .S0 (nx36179)) ;
    mux21_ni ix14797 (.Y (nx14796), .A0 (mdr_data_out[7]), .A1 (
             booth_booth_integration_output_7_8), .S0 (nx36189)) ;
    mux21_ni ix22974 (.Y (nx22973), .A0 (booth_booth_integration_output_7_8), .A1 (
             nx14784), .S0 (nx36179)) ;
    mux21_ni ix14785 (.Y (nx14784), .A0 (mdr_data_out[8]), .A1 (
             booth_booth_integration_output_7_9), .S0 (nx36189)) ;
    mux21_ni ix22964 (.Y (nx22963), .A0 (booth_booth_integration_output_7_9), .A1 (
             nx14772), .S0 (nx36179)) ;
    mux21_ni ix14773 (.Y (nx14772), .A0 (mdr_data_out[9]), .A1 (
             booth_booth_integration_output_7_10), .S0 (nx36189)) ;
    mux21_ni ix22954 (.Y (nx22953), .A0 (booth_booth_integration_output_7_10), .A1 (
             nx14760), .S0 (nx36181)) ;
    mux21_ni ix14761 (.Y (nx14760), .A0 (mdr_data_out[10]), .A1 (
             booth_booth_integration_output_7_11), .S0 (nx36189)) ;
    mux21_ni ix22944 (.Y (nx22943), .A0 (booth_booth_integration_output_7_11), .A1 (
             nx14748), .S0 (nx36181)) ;
    mux21_ni ix14749 (.Y (nx14748), .A0 (mdr_data_out[11]), .A1 (
             booth_booth_integration_output_7_12), .S0 (nx36189)) ;
    mux21_ni ix22934 (.Y (nx22933), .A0 (booth_booth_integration_output_7_12), .A1 (
             nx14736), .S0 (nx36181)) ;
    mux21_ni ix14737 (.Y (nx14736), .A0 (mdr_data_out[12]), .A1 (
             booth_booth_integration_output_7_13), .S0 (nx36191)) ;
    mux21_ni ix22924 (.Y (nx22923), .A0 (booth_booth_integration_output_7_13), .A1 (
             nx14724), .S0 (nx36181)) ;
    mux21_ni ix14725 (.Y (nx14724), .A0 (mdr_data_out[13]), .A1 (
             booth_booth_integration_output_7_14), .S0 (nx36191)) ;
    mux21_ni ix22914 (.Y (nx22913), .A0 (booth_booth_integration_output_7_14), .A1 (
             nx14712), .S0 (nx36181)) ;
    mux21_ni ix14713 (.Y (nx14712), .A0 (mdr_data_out[14]), .A1 (
             booth_booth_integration_output_7_15), .S0 (nx36191)) ;
    mux21 ix22904 (.Y (nx22903), .A0 (nx31848), .A1 (nx31490), .S0 (nx36181)) ;
    mux21_ni ix22554 (.Y (nx22553), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_0), .A1 (nx35043), .S0 (
             nx35839)) ;
    and02 ix22540 (.Y (nx22539), .A0 (nx36361), .A1 (
          booth_booth_integrtaion_7_shift_Reg_count_0)) ;
    mux21_ni ix22734 (.Y (nx22733), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_9), .A1 (nx35029), .S0 (
             nx35839)) ;
    mux21_ni ix22724 (.Y (nx22723), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_9), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_8), .S0 (nx36181)) ;
    mux21_ni ix22714 (.Y (nx22713), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_8), .S0 (nx35839)) ;
    mux21_ni ix22704 (.Y (nx22703), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_8), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_7), .S0 (nx36183)) ;
    mux21_ni ix22694 (.Y (nx22693), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_7), .S0 (nx35839)) ;
    mux21_ni ix22684 (.Y (nx22683), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_7), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_6), .S0 (nx36183)) ;
    mux21_ni ix22674 (.Y (nx22673), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_6), .S0 (nx35839)) ;
    mux21_ni ix22664 (.Y (nx22663), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_6), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_5), .S0 (nx36183)) ;
    mux21_ni ix22654 (.Y (nx22653), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_5), .S0 (nx35839)) ;
    mux21_ni ix22644 (.Y (nx22643), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_5), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_4), .S0 (nx36183)) ;
    mux21_ni ix22634 (.Y (nx22633), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_4), .S0 (nx35841)) ;
    mux21_ni ix22624 (.Y (nx22623), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_4), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_3), .S0 (nx36183)) ;
    mux21_ni ix22614 (.Y (nx22613), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_3), .S0 (nx35841)) ;
    mux21_ni ix22604 (.Y (nx22603), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_3), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_2), .S0 (nx36183)) ;
    mux21_ni ix22594 (.Y (nx22593), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_2), .S0 (nx35841)) ;
    mux21_ni ix22584 (.Y (nx22583), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_2), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_1), .S0 (nx36183)) ;
    mux21_ni ix22574 (.Y (nx22573), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_1), .A1 (
             booth_booth_integrtaion_7_shift_Reg_output_1), .S0 (nx35841)) ;
    mux21_ni ix22564 (.Y (nx22563), .A0 (
             booth_booth_integrtaion_7_shift_Reg_count_1), .A1 (nx35043), .S0 (
             nx36185)) ;
    and02 ix14153 (.Y (nx14152), .A0 (nx31563), .A1 (nx35775)) ;
    or03 ix31566 (.Y (nx31565), .A0 (nx31567), .A1 (
         booth_booth_integrtaion_7_shift_reg_output_0), .A2 (nx36361)) ;
    mux21_ni ix22894 (.Y (nx22893), .A0 (
             booth_booth_integrtaion_7_booth_output_16), .A1 (nx14682), .S0 (
             nx36185)) ;
    nor02ii ix14683 (.Y (nx14682), .A0 (nx31574), .A1 (nx36191)) ;
    nor02ii ix14159 (.Y (nx14158), .A0 (nx31558), .A1 (
            booth_booth_integrtaion_7_booth_output_16)) ;
    xor2 ix14677 (.Y (nx13334), .A0 (nx31580), .A1 (nx31844)) ;
    xor2 ix14665 (.Y (nx13335), .A0 (nx31605), .A1 (nx35563)) ;
    mux21_ni ix22874 (.Y (nx22873), .A0 (
             booth_booth_integrtaion_7_booth_output_18), .A1 (nx14658), .S0 (
             nx36185)) ;
    nor02ii ix14659 (.Y (nx14658), .A0 (nx31595), .A1 (nx36191)) ;
    xor2 ix14653 (.Y (nx13336), .A0 (nx31610), .A1 (nx31841)) ;
    or02 ix31627 (.Y (nx31626), .A0 (nx31563), .A1 (nx35777)) ;
    xor2 ix14641 (.Y (nx13337), .A0 (nx31644), .A1 (nx35565)) ;
    mux21_ni ix22854 (.Y (nx22853), .A0 (
             booth_booth_integrtaion_7_booth_output_20), .A1 (nx14634), .S0 (
             nx36185)) ;
    nor02ii ix14635 (.Y (nx14634), .A0 (nx31632), .A1 (nx36191)) ;
    xor2 ix14629 (.Y (nx13339), .A0 (nx31649), .A1 (nx31838)) ;
    xor2 ix14617 (.Y (nx13341), .A0 (nx31679), .A1 (nx35567)) ;
    mux21_ni ix22834 (.Y (nx22833), .A0 (
             booth_booth_integrtaion_7_booth_output_22), .A1 (nx14610), .S0 (
             nx36185)) ;
    nor02ii ix14611 (.Y (nx14610), .A0 (nx31667), .A1 (nx36191)) ;
    xor2 ix14605 (.Y (nx13343), .A0 (nx31684), .A1 (nx31835)) ;
    xor2 ix14593 (.Y (nx13344), .A0 (nx31714), .A1 (nx35569)) ;
    mux21_ni ix22814 (.Y (nx22813), .A0 (
             booth_booth_integrtaion_7_booth_output_24), .A1 (nx14586), .S0 (
             nx36185)) ;
    nor02ii ix14587 (.Y (nx14586), .A0 (nx31702), .A1 (nx36193)) ;
    xor2 ix14581 (.Y (nx13345), .A0 (nx31719), .A1 (nx31832)) ;
    xor2 ix14569 (.Y (nx13346), .A0 (nx31749), .A1 (nx35571)) ;
    mux21_ni ix22794 (.Y (nx22793), .A0 (
             booth_booth_integrtaion_7_booth_output_26), .A1 (nx14562), .S0 (
             nx36185)) ;
    nor02ii ix14563 (.Y (nx14562), .A0 (nx31737), .A1 (nx36193)) ;
    xor2 ix14557 (.Y (nx13347), .A0 (nx31754), .A1 (nx31829)) ;
    xor2 ix14545 (.Y (nx13348), .A0 (nx31784), .A1 (nx35573)) ;
    mux21_ni ix22774 (.Y (nx22773), .A0 (
             booth_booth_integrtaion_7_booth_output_28), .A1 (nx14538), .S0 (
             nx35555)) ;
    nor02ii ix14539 (.Y (nx14538), .A0 (nx31772), .A1 (nx36193)) ;
    xor2 ix14533 (.Y (nx13349), .A0 (nx31789), .A1 (nx31826)) ;
    xor2 ix14521 (.Y (nx13351), .A0 (nx31819), .A1 (nx35575)) ;
    mux21_ni ix22754 (.Y (nx22753), .A0 (
             booth_booth_integrtaion_7_booth_output_31), .A1 (nx14514), .S0 (
             nx35555)) ;
    nor02ii ix14515 (.Y (nx14514), .A0 (nx31807), .A1 (nx36193)) ;
    xor2 ix14509 (.Y (nx14508), .A0 (nx31819), .A1 (nx31822)) ;
    nor02ii ix14695 (.Y (nx14694), .A0 (nx14158), .A1 (nx36193)) ;
    or03 ix31873 (.Y (nx31872), .A0 (nx32056), .A1 (nx36199), .A2 (nx36073)) ;
    mux21_ni ix23344 (.Y (nx23343), .A0 (label_8_output[14]), .A1 (
             label_8_input_14), .S0 (nx36259)) ;
    mux21_ni ix15339 (.Y (nx15338), .A0 (nx15334), .A1 (
             label_8_input_state_machine_14), .S0 (nx35937)) ;
    mux21_ni ix22524 (.Y (nx22523), .A0 (label_8_input_state_machine_14), .A1 (
             mdr_data_out[126]), .S0 (nx36221)) ;
    mux21_ni ix23334 (.Y (nx23333), .A0 (label_8_output[13]), .A1 (
             label_8_input_13), .S0 (nx36259)) ;
    mux21_ni ix15313 (.Y (nx15312), .A0 (nx15308), .A1 (
             label_8_input_state_machine_13), .S0 (nx35937)) ;
    mux21_ni ix23324 (.Y (nx23323), .A0 (label_8_input_state_machine_13), .A1 (
             mdr_data_out[125]), .S0 (nx36221)) ;
    mux21_ni ix23294 (.Y (nx23293), .A0 (label_8_output[11]), .A1 (
             label_8_input_11), .S0 (nx36259)) ;
    mux21_ni ix15249 (.Y (nx15248), .A0 (nx15244), .A1 (
             label_8_input_state_machine_11), .S0 (nx35937)) ;
    mux21_ni ix23284 (.Y (nx23283), .A0 (label_8_input_state_machine_11), .A1 (
             mdr_data_out[123]), .S0 (nx36221)) ;
    mux21_ni ix23254 (.Y (nx23253), .A0 (label_8_output[9]), .A1 (
             label_8_input_9), .S0 (nx36259)) ;
    mux21_ni ix15185 (.Y (nx15184), .A0 (nx15180), .A1 (
             label_8_input_state_machine_9), .S0 (nx35937)) ;
    mux21_ni ix23244 (.Y (nx23243), .A0 (label_8_input_state_machine_9), .A1 (
             mdr_data_out[121]), .S0 (nx36221)) ;
    mux21_ni ix23214 (.Y (nx23213), .A0 (label_8_output[7]), .A1 (
             label_8_input_7), .S0 (nx36259)) ;
    mux21_ni ix15121 (.Y (nx15120), .A0 (nx15116), .A1 (
             label_8_input_state_machine_7), .S0 (nx35937)) ;
    mux21_ni ix23204 (.Y (nx23203), .A0 (label_8_input_state_machine_7), .A1 (
             mdr_data_out[119]), .S0 (nx36221)) ;
    mux21_ni ix23174 (.Y (nx23173), .A0 (label_8_output[5]), .A1 (
             label_8_input_5), .S0 (nx36259)) ;
    mux21_ni ix15057 (.Y (nx15056), .A0 (nx15052), .A1 (
             label_8_input_state_machine_5), .S0 (nx35937)) ;
    mux21_ni ix23164 (.Y (nx23163), .A0 (label_8_input_state_machine_5), .A1 (
             mdr_data_out[117]), .S0 (nx36221)) ;
    mux21_ni ix23134 (.Y (nx23133), .A0 (label_8_output[3]), .A1 (
             label_8_input_3), .S0 (nx36259)) ;
    mux21_ni ix14993 (.Y (nx14992), .A0 (nx14988), .A1 (
             label_8_input_state_machine_3), .S0 (nx35935)) ;
    mux21_ni ix23124 (.Y (nx23123), .A0 (label_8_input_state_machine_3), .A1 (
             mdr_data_out[115]), .S0 (nx36223)) ;
    mux21_ni ix23094 (.Y (nx23093), .A0 (label_8_output[1]), .A1 (
             label_8_input_1), .S0 (nx36261)) ;
    mux21_ni ix14929 (.Y (nx14928), .A0 (nx14924), .A1 (
             label_8_input_state_machine_1), .S0 (nx35935)) ;
    mux21_ni ix23084 (.Y (nx23083), .A0 (label_8_input_state_machine_1), .A1 (
             mdr_data_out[113]), .S0 (nx36223)) ;
    xnor2 ix31965 (.Y (nx31964), .A0 (nx31862), .A1 (nx31974)) ;
    mux21_ni ix23114 (.Y (nx23113), .A0 (label_8_output[2]), .A1 (
             label_8_input_2), .S0 (nx36261)) ;
    mux21_ni ix14961 (.Y (nx14960), .A0 (nx14956), .A1 (
             label_8_input_state_machine_2), .S0 (nx35167)) ;
    mux21_ni ix23104 (.Y (nx23103), .A0 (label_8_input_state_machine_2), .A1 (
             mdr_data_out[114]), .S0 (nx36223)) ;
    xnor2 ix31980 (.Y (nx31979), .A0 (nx31860), .A1 (nx31989)) ;
    mux21_ni ix23154 (.Y (nx23153), .A0 (label_8_output[4]), .A1 (
             label_8_input_4), .S0 (nx36261)) ;
    mux21_ni ix15025 (.Y (nx15024), .A0 (nx15020), .A1 (
             label_8_input_state_machine_4), .S0 (nx35167)) ;
    mux21_ni ix23144 (.Y (nx23143), .A0 (label_8_input_state_machine_4), .A1 (
             mdr_data_out[116]), .S0 (nx36223)) ;
    xnor2 ix31995 (.Y (nx31994), .A0 (nx31858), .A1 (nx32004)) ;
    mux21_ni ix23194 (.Y (nx23193), .A0 (label_8_output[6]), .A1 (
             label_8_input_6), .S0 (nx36261)) ;
    mux21_ni ix15089 (.Y (nx15088), .A0 (nx15084), .A1 (
             label_8_input_state_machine_6), .S0 (nx35937)) ;
    mux21_ni ix23184 (.Y (nx23183), .A0 (label_8_input_state_machine_6), .A1 (
             mdr_data_out[118]), .S0 (nx36223)) ;
    xnor2 ix32010 (.Y (nx32009), .A0 (nx31856), .A1 (nx32019)) ;
    mux21_ni ix23234 (.Y (nx23233), .A0 (label_8_output[8]), .A1 (
             label_8_input_8), .S0 (nx36261)) ;
    mux21_ni ix15153 (.Y (nx15152), .A0 (nx15148), .A1 (
             label_8_input_state_machine_8), .S0 (nx35939)) ;
    mux21_ni ix23224 (.Y (nx23223), .A0 (label_8_input_state_machine_8), .A1 (
             mdr_data_out[120]), .S0 (nx36223)) ;
    xnor2 ix32025 (.Y (nx32024), .A0 (nx31854), .A1 (nx32034)) ;
    mux21_ni ix23274 (.Y (nx23273), .A0 (label_8_output[10]), .A1 (
             label_8_input_10), .S0 (nx36261)) ;
    mux21_ni ix15217 (.Y (nx15216), .A0 (nx15212), .A1 (
             label_8_input_state_machine_10), .S0 (nx35939)) ;
    mux21_ni ix23264 (.Y (nx23263), .A0 (label_8_input_state_machine_10), .A1 (
             mdr_data_out[122]), .S0 (nx36223)) ;
    xnor2 ix32040 (.Y (nx32039), .A0 (nx31852), .A1 (nx32049)) ;
    mux21_ni ix23314 (.Y (nx23313), .A0 (label_8_output[12]), .A1 (
             label_8_input_12), .S0 (nx36261)) ;
    mux21_ni ix15281 (.Y (nx15280), .A0 (nx15276), .A1 (
             label_8_input_state_machine_12), .S0 (nx35939)) ;
    mux21_ni ix23304 (.Y (nx23303), .A0 (label_8_input_state_machine_12), .A1 (
             mdr_data_out[124]), .S0 (nx35597)) ;
    xnor2 ix32055 (.Y (nx32054), .A0 (nx31850), .A1 (nx32056)) ;
    or03 ix32062 (.Y (nx32061), .A0 (nx32245), .A1 (nx36125), .A2 (nx36073)) ;
    mux21_ni ix22504 (.Y (nx22503), .A0 (label_7_output[14]), .A1 (
             label_7_input_14), .S0 (nx36263)) ;
    mux21_ni ix14023 (.Y (nx14022), .A0 (nx14018), .A1 (
             label_7_input_state_machine_14), .S0 (nx35939)) ;
    mux21_ni ix21684 (.Y (nx21683), .A0 (label_7_input_state_machine_14), .A1 (
             mdr_data_out[110]), .S0 (nx35597)) ;
    mux21_ni ix22494 (.Y (nx22493), .A0 (label_7_output[13]), .A1 (
             label_7_input_13), .S0 (nx36263)) ;
    mux21_ni ix13997 (.Y (nx13996), .A0 (nx13992), .A1 (
             label_7_input_state_machine_13), .S0 (nx35939)) ;
    mux21_ni ix22484 (.Y (nx22483), .A0 (label_7_input_state_machine_13), .A1 (
             mdr_data_out[109]), .S0 (nx35597)) ;
    mux21_ni ix22454 (.Y (nx22453), .A0 (label_7_output[11]), .A1 (
             label_7_input_11), .S0 (nx36263)) ;
    mux21_ni ix13933 (.Y (nx13932), .A0 (nx13928), .A1 (
             label_7_input_state_machine_11), .S0 (nx35939)) ;
    mux21_ni ix22444 (.Y (nx22443), .A0 (label_7_input_state_machine_11), .A1 (
             mdr_data_out[107]), .S0 (nx35597)) ;
    mux21_ni ix22414 (.Y (nx22413), .A0 (label_7_output[9]), .A1 (
             label_7_input_9), .S0 (nx36263)) ;
    mux21_ni ix13869 (.Y (nx13868), .A0 (nx13864), .A1 (
             label_7_input_state_machine_9), .S0 (nx35939)) ;
    mux21_ni ix22404 (.Y (nx22403), .A0 (label_7_input_state_machine_9), .A1 (
             mdr_data_out[105]), .S0 (nx35597)) ;
    mux21_ni ix22374 (.Y (nx22373), .A0 (label_7_output[7]), .A1 (
             label_7_input_7), .S0 (nx36263)) ;
    mux21_ni ix13805 (.Y (nx13804), .A0 (nx13800), .A1 (
             label_7_input_state_machine_7), .S0 (nx35941)) ;
    mux21_ni ix22364 (.Y (nx22363), .A0 (label_7_input_state_machine_7), .A1 (
             mdr_data_out[103]), .S0 (nx35597)) ;
    mux21_ni ix22334 (.Y (nx22333), .A0 (label_7_output[5]), .A1 (
             label_7_input_5), .S0 (nx36263)) ;
    mux21_ni ix13741 (.Y (nx13740), .A0 (nx13736), .A1 (
             label_7_input_state_machine_5), .S0 (nx35941)) ;
    mux21_ni ix22324 (.Y (nx22323), .A0 (label_7_input_state_machine_5), .A1 (
             mdr_data_out[101]), .S0 (nx35597)) ;
    mux21_ni ix22294 (.Y (nx22293), .A0 (label_7_output[3]), .A1 (
             label_7_input_3), .S0 (nx36263)) ;
    mux21_ni ix13677 (.Y (nx13676), .A0 (nx13672), .A1 (
             label_7_input_state_machine_3), .S0 (nx35941)) ;
    mux21_ni ix22284 (.Y (nx22283), .A0 (label_7_input_state_machine_3), .A1 (
             mdr_data_out[99]), .S0 (nx36225)) ;
    mux21_ni ix22254 (.Y (nx22253), .A0 (label_7_output[1]), .A1 (
             label_7_input_1), .S0 (nx35605)) ;
    mux21_ni ix13613 (.Y (nx13612), .A0 (nx13608), .A1 (
             label_7_input_state_machine_1), .S0 (nx35941)) ;
    mux21_ni ix22244 (.Y (nx22243), .A0 (label_7_input_state_machine_1), .A1 (
             mdr_data_out[97]), .S0 (nx36225)) ;
    xnor2 ix32154 (.Y (nx32153), .A0 (nx31423), .A1 (nx32163)) ;
    mux21_ni ix22274 (.Y (nx22273), .A0 (label_7_output[2]), .A1 (
             label_7_input_2), .S0 (nx35605)) ;
    mux21_ni ix13645 (.Y (nx13644), .A0 (nx13640), .A1 (
             label_7_input_state_machine_2), .S0 (nx35941)) ;
    mux21_ni ix22264 (.Y (nx22263), .A0 (label_7_input_state_machine_2), .A1 (
             mdr_data_out[98]), .S0 (nx36225)) ;
    xnor2 ix32169 (.Y (nx32168), .A0 (nx31421), .A1 (nx32178)) ;
    mux21_ni ix22314 (.Y (nx22313), .A0 (label_7_output[4]), .A1 (
             label_7_input_4), .S0 (nx35605)) ;
    mux21_ni ix13709 (.Y (nx13708), .A0 (nx13704), .A1 (
             label_7_input_state_machine_4), .S0 (nx35941)) ;
    mux21_ni ix22304 (.Y (nx22303), .A0 (label_7_input_state_machine_4), .A1 (
             mdr_data_out[100]), .S0 (nx36225)) ;
    xnor2 ix32184 (.Y (nx32183), .A0 (nx31419), .A1 (nx32193)) ;
    mux21_ni ix22354 (.Y (nx22353), .A0 (label_7_output[6]), .A1 (
             label_7_input_6), .S0 (nx35605)) ;
    mux21_ni ix13773 (.Y (nx13772), .A0 (nx13768), .A1 (
             label_7_input_state_machine_6), .S0 (nx35941)) ;
    mux21_ni ix22344 (.Y (nx22343), .A0 (label_7_input_state_machine_6), .A1 (
             mdr_data_out[102]), .S0 (nx36225)) ;
    xnor2 ix32199 (.Y (nx32198), .A0 (nx31417), .A1 (nx32208)) ;
    mux21_ni ix22394 (.Y (nx22393), .A0 (label_7_output[8]), .A1 (
             label_7_input_8), .S0 (nx35605)) ;
    mux21_ni ix13837 (.Y (nx13836), .A0 (nx13832), .A1 (
             label_7_input_state_machine_8), .S0 (nx35943)) ;
    mux21_ni ix22384 (.Y (nx22383), .A0 (label_7_input_state_machine_8), .A1 (
             mdr_data_out[104]), .S0 (nx36225)) ;
    xnor2 ix32214 (.Y (nx32213), .A0 (nx31415), .A1 (nx32223)) ;
    mux21_ni ix22434 (.Y (nx22433), .A0 (label_7_output[10]), .A1 (
             label_7_input_10), .S0 (nx35605)) ;
    mux21_ni ix13901 (.Y (nx13900), .A0 (nx13896), .A1 (
             label_7_input_state_machine_10), .S0 (nx35943)) ;
    mux21_ni ix22424 (.Y (nx22423), .A0 (label_7_input_state_machine_10), .A1 (
             mdr_data_out[106]), .S0 (nx36225)) ;
    xnor2 ix32229 (.Y (nx32228), .A0 (nx31413), .A1 (nx32238)) ;
    mux21_ni ix22474 (.Y (nx22473), .A0 (label_7_output[12]), .A1 (
             label_7_input_12), .S0 (nx35605)) ;
    mux21_ni ix13965 (.Y (nx13964), .A0 (nx13960), .A1 (
             label_7_input_state_machine_12), .S0 (nx35943)) ;
    mux21_ni ix22464 (.Y (nx22463), .A0 (label_7_input_state_machine_12), .A1 (
             mdr_data_out[108]), .S0 (nx36227)) ;
    xnor2 ix32244 (.Y (nx32243), .A0 (nx31411), .A1 (nx32245)) ;
    xnor2 ix15361 (.Y (nx15360), .A0 (nx31869), .A1 (nx32059)) ;
    xnor2 ix32249 (.Y (nx32248), .A0 (nx32252), .A1 (
          max_calc_comparator_fourth_inp1_13)) ;
    or03 ix32267 (.Y (nx32266), .A0 (nx32049), .A1 (nx36125), .A2 (nx36073)) ;
    or03 ix32273 (.Y (nx32272), .A0 (nx32238), .A1 (nx36125), .A2 (nx36073)) ;
    xnor2 ix15405 (.Y (nx15404), .A0 (nx32263), .A1 (nx32270)) ;
    xnor2 ix32277 (.Y (nx32276), .A0 (nx32280), .A1 (
          max_calc_comparator_fourth_inp1_11)) ;
    or03 ix32295 (.Y (nx32294), .A0 (nx32034), .A1 (nx36127), .A2 (nx36073)) ;
    or03 ix32301 (.Y (nx32300), .A0 (nx32223), .A1 (nx36127), .A2 (nx36073)) ;
    xnor2 ix15449 (.Y (nx15448), .A0 (nx32291), .A1 (nx32298)) ;
    xnor2 ix32305 (.Y (nx32304), .A0 (nx32308), .A1 (
          max_calc_comparator_fourth_inp1_9)) ;
    or03 ix32323 (.Y (nx32322), .A0 (nx32019), .A1 (nx36127), .A2 (nx35367)) ;
    or03 ix32329 (.Y (nx32328), .A0 (nx32208), .A1 (nx36127), .A2 (nx35367)) ;
    xnor2 ix15493 (.Y (nx15492), .A0 (nx32319), .A1 (nx32326)) ;
    xnor2 ix32333 (.Y (nx32332), .A0 (nx32336), .A1 (
          max_calc_comparator_fourth_inp1_7)) ;
    or03 ix32351 (.Y (nx32350), .A0 (nx32004), .A1 (nx36127), .A2 (nx35369)) ;
    or03 ix32357 (.Y (nx32356), .A0 (nx32193), .A1 (nx36127), .A2 (nx35369)) ;
    xnor2 ix15537 (.Y (nx15536), .A0 (nx32347), .A1 (nx32354)) ;
    xnor2 ix32361 (.Y (nx32360), .A0 (nx32364), .A1 (
          max_calc_comparator_fourth_inp1_5)) ;
    or03 ix32379 (.Y (nx32378), .A0 (nx31989), .A1 (nx36127), .A2 (nx35369)) ;
    or03 ix32385 (.Y (nx32384), .A0 (nx32178), .A1 (nx36129), .A2 (nx35369)) ;
    xnor2 ix15581 (.Y (nx15580), .A0 (nx32375), .A1 (nx32382)) ;
    xnor2 ix32389 (.Y (nx32388), .A0 (nx32392), .A1 (
          max_calc_comparator_fourth_inp1_3)) ;
    or03 ix32407 (.Y (nx32406), .A0 (nx31974), .A1 (nx36129), .A2 (nx35369)) ;
    or03 ix32413 (.Y (nx32412), .A0 (nx32163), .A1 (nx36129), .A2 (nx35369)) ;
    xnor2 ix15625 (.Y (nx15624), .A0 (nx32403), .A1 (nx32410)) ;
    xnor2 ix15647 (.Y (nx15646), .A0 (nx32418), .A1 (nx32422)) ;
    xnor2 ix15873 (.Y (nx15872), .A0 (nx32433), .A1 (nx32451)) ;
    mux21_ni ix23654 (.Y (nx23653), .A0 (label_8_output[15]), .A1 (
             label_8_input_15), .S0 (nx36265)) ;
    mux21_ni ix15809 (.Y (nx15808), .A0 (nx15804), .A1 (
             label_8_input_state_machine_15), .S0 (nx35943)) ;
    mux21_ni ix23644 (.Y (nx23643), .A0 (label_8_input_state_machine_15), .A1 (
             mdr_data_out[127]), .S0 (nx36227)) ;
    xor2 ix32447 (.Y (nx32446), .A0 (nx31848), .A1 (label_8_output[15])) ;
    or03 ix32454 (.Y (nx32453), .A0 (nx35649), .A1 (nx36129), .A2 (nx35369)) ;
    inv01 ix35648 (.Y (nx35649), .A (label_7_output[15])) ;
    mux21_ni ix23684 (.Y (nx23683), .A0 (label_7_output[15]), .A1 (
             label_7_input_15), .S0 (nx36265)) ;
    mux21_ni ix15851 (.Y (nx15850), .A0 (nx15846), .A1 (
             label_7_input_state_machine_15), .S0 (nx35943)) ;
    mux21_ni ix23674 (.Y (nx23673), .A0 (label_7_input_state_machine_15), .A1 (
             mdr_data_out[111]), .S0 (nx36227)) ;
    xor2 ix32465 (.Y (nx32464), .A0 (nx31409), .A1 (label_7_output[15])) ;
    mux21 ix15897 (.Y (nx15896), .A0 (nx32665), .A1 (nx32660), .S0 (nx35979)) ;
    mux21_ni ix14954 (.Y (nx14953), .A0 (label_4_output[14]), .A1 (
             label_4_input_14), .S0 (nx36265)) ;
    mux21_ni ix2187 (.Y (nx2186), .A0 (nx2182), .A1 (
             label_4_input_state_machine_14), .S0 (nx35943)) ;
    mux21_ni ix14944 (.Y (nx14943), .A0 (label_4_input_state_machine_14), .A1 (
             mdr_data_out[62]), .S0 (nx36227)) ;
    mux21_ni ix14934 (.Y (nx14933), .A0 (label_4_output[13]), .A1 (
             label_4_input_13), .S0 (nx36265)) ;
    mux21_ni ix2155 (.Y (nx2154), .A0 (nx2150), .A1 (
             label_4_input_state_machine_13), .S0 (nx35943)) ;
    mux21_ni ix14924 (.Y (nx14923), .A0 (label_4_input_state_machine_13), .A1 (
             mdr_data_out[61]), .S0 (nx36227)) ;
    mux21_ni ix14894 (.Y (nx14893), .A0 (label_4_output[11]), .A1 (
             label_4_input_11), .S0 (nx36265)) ;
    mux21_ni ix2091 (.Y (nx2090), .A0 (nx2086), .A1 (
             label_4_input_state_machine_11), .S0 (nx35945)) ;
    mux21_ni ix14884 (.Y (nx14883), .A0 (label_4_input_state_machine_11), .A1 (
             mdr_data_out[59]), .S0 (nx36227)) ;
    mux21_ni ix14854 (.Y (nx14853), .A0 (label_4_output[9]), .A1 (
             label_4_input_9), .S0 (nx36265)) ;
    mux21_ni ix2027 (.Y (nx2026), .A0 (nx2022), .A1 (
             label_4_input_state_machine_9), .S0 (nx35945)) ;
    mux21_ni ix14844 (.Y (nx14843), .A0 (label_4_input_state_machine_9), .A1 (
             mdr_data_out[57]), .S0 (nx36227)) ;
    mux21_ni ix14814 (.Y (nx14813), .A0 (label_4_output[7]), .A1 (
             label_4_input_7), .S0 (nx36265)) ;
    mux21_ni ix1963 (.Y (nx1962), .A0 (nx1958), .A1 (
             label_4_input_state_machine_7), .S0 (nx35945)) ;
    mux21_ni ix14804 (.Y (nx14803), .A0 (label_4_input_state_machine_7), .A1 (
             mdr_data_out[55]), .S0 (nx36229)) ;
    mux21_ni ix14774 (.Y (nx14773), .A0 (label_4_output[5]), .A1 (
             label_4_input_5), .S0 (nx36267)) ;
    mux21_ni ix1899 (.Y (nx1898), .A0 (nx1894), .A1 (
             label_4_input_state_machine_5), .S0 (nx35945)) ;
    mux21_ni ix14764 (.Y (nx14763), .A0 (label_4_input_state_machine_5), .A1 (
             mdr_data_out[53]), .S0 (nx36229)) ;
    mux21_ni ix14734 (.Y (nx14733), .A0 (label_4_output[3]), .A1 (
             label_4_input_3), .S0 (nx36267)) ;
    mux21_ni ix1835 (.Y (nx1834), .A0 (nx1830), .A1 (
             label_4_input_state_machine_3), .S0 (nx35945)) ;
    mux21_ni ix14724 (.Y (nx14723), .A0 (label_4_input_state_machine_3), .A1 (
             mdr_data_out[51]), .S0 (nx36229)) ;
    mux21_ni ix14694 (.Y (nx14693), .A0 (label_4_output[1]), .A1 (
             label_4_input_1), .S0 (nx36267)) ;
    mux21_ni ix1771 (.Y (nx1770), .A0 (nx1766), .A1 (
             label_4_input_state_machine_1), .S0 (nx35945)) ;
    mux21_ni ix14684 (.Y (nx14683), .A0 (label_4_input_state_machine_1), .A1 (
             mdr_data_out[49]), .S0 (nx36229)) ;
    xnor2 ix32569 (.Y (nx32568), .A0 (nx30980), .A1 (nx32578)) ;
    mux21_ni ix14714 (.Y (nx14713), .A0 (label_4_output[2]), .A1 (
             label_4_input_2), .S0 (nx36267)) ;
    mux21_ni ix1803 (.Y (nx1802), .A0 (nx1798), .A1 (
             label_4_input_state_machine_2), .S0 (nx35945)) ;
    mux21_ni ix14704 (.Y (nx14703), .A0 (label_4_input_state_machine_2), .A1 (
             mdr_data_out[50]), .S0 (nx36229)) ;
    xnor2 ix32584 (.Y (nx32583), .A0 (nx30978), .A1 (nx32593)) ;
    mux21_ni ix14754 (.Y (nx14753), .A0 (label_4_output[4]), .A1 (
             label_4_input_4), .S0 (nx36267)) ;
    mux21_ni ix1867 (.Y (nx1866), .A0 (nx1862), .A1 (
             label_4_input_state_machine_4), .S0 (nx35947)) ;
    mux21_ni ix14744 (.Y (nx14743), .A0 (label_4_input_state_machine_4), .A1 (
             mdr_data_out[52]), .S0 (nx36229)) ;
    xnor2 ix32599 (.Y (nx32598), .A0 (nx30976), .A1 (nx32608)) ;
    mux21_ni ix14794 (.Y (nx14793), .A0 (label_4_output[6]), .A1 (
             label_4_input_6), .S0 (nx36267)) ;
    mux21_ni ix1931 (.Y (nx1930), .A0 (nx1926), .A1 (
             label_4_input_state_machine_6), .S0 (nx35947)) ;
    mux21_ni ix14784 (.Y (nx14783), .A0 (label_4_input_state_machine_6), .A1 (
             mdr_data_out[54]), .S0 (nx36229)) ;
    xnor2 ix32614 (.Y (nx32613), .A0 (nx30974), .A1 (nx32623)) ;
    mux21_ni ix14834 (.Y (nx14833), .A0 (label_4_output[8]), .A1 (
             label_4_input_8), .S0 (nx36267)) ;
    mux21_ni ix1995 (.Y (nx1994), .A0 (nx1990), .A1 (
             label_4_input_state_machine_8), .S0 (nx35947)) ;
    mux21_ni ix14824 (.Y (nx14823), .A0 (label_4_input_state_machine_8), .A1 (
             mdr_data_out[56]), .S0 (nx36231)) ;
    xnor2 ix32629 (.Y (nx32628), .A0 (nx30972), .A1 (nx32638)) ;
    mux21_ni ix14874 (.Y (nx14873), .A0 (label_4_output[10]), .A1 (
             label_4_input_10), .S0 (nx36269)) ;
    mux21_ni ix2059 (.Y (nx2058), .A0 (nx2054), .A1 (
             label_4_input_state_machine_10), .S0 (nx35947)) ;
    mux21_ni ix14864 (.Y (nx14863), .A0 (label_4_input_state_machine_10), .A1 (
             mdr_data_out[58]), .S0 (nx36231)) ;
    xnor2 ix32644 (.Y (nx32643), .A0 (nx30970), .A1 (nx32653)) ;
    mux21_ni ix14914 (.Y (nx14913), .A0 (label_4_output[12]), .A1 (
             label_4_input_12), .S0 (nx36269)) ;
    mux21_ni ix2123 (.Y (nx2122), .A0 (nx2118), .A1 (
             label_4_input_state_machine_12), .S0 (nx35947)) ;
    mux21_ni ix14904 (.Y (nx14903), .A0 (label_4_input_state_machine_12), .A1 (
             mdr_data_out[60]), .S0 (nx36231)) ;
    xnor2 ix32659 (.Y (nx32658), .A0 (nx30968), .A1 (nx32660)) ;
    ao32 ix23704 (.Y (nx23703), .A0 (nx35961), .A1 (nx35651), .A2 (nx36291), .B0 (
         max_calc_ans4_14), .B1 (nx35877)) ;
    mux21 ix32664 (.Y (nx35651), .A0 (nx31869), .A1 (nx32059), .S0 (nx35893)) ;
    mux21 ix12713 (.Y (nx12712), .A0 (nx32861), .A1 (nx32856), .S0 (nx35979)) ;
    mux21_ni ix15804 (.Y (nx15803), .A0 (label_3_output[14]), .A1 (
             label_3_input_14), .S0 (nx36269)) ;
    mux21_ni ix3525 (.Y (nx3524), .A0 (nx3520), .A1 (
             label_3_input_state_machine_14), .S0 (nx35949)) ;
    mux21_ni ix15794 (.Y (nx15793), .A0 (label_3_input_state_machine_14), .A1 (
             mdr_data_out[46]), .S0 (nx36231)) ;
    mux21_ni ix15784 (.Y (nx15783), .A0 (label_3_output[13]), .A1 (
             label_3_input_13), .S0 (nx36269)) ;
    mux21_ni ix3493 (.Y (nx3492), .A0 (nx3488), .A1 (
             label_3_input_state_machine_13), .S0 (nx35949)) ;
    mux21_ni ix15774 (.Y (nx15773), .A0 (label_3_input_state_machine_13), .A1 (
             mdr_data_out[45]), .S0 (nx36231)) ;
    mux21_ni ix15744 (.Y (nx15743), .A0 (label_3_output[11]), .A1 (
             label_3_input_11), .S0 (nx36269)) ;
    mux21_ni ix3429 (.Y (nx3428), .A0 (nx3424), .A1 (
             label_3_input_state_machine_11), .S0 (nx35949)) ;
    mux21_ni ix15734 (.Y (nx15733), .A0 (label_3_input_state_machine_11), .A1 (
             mdr_data_out[43]), .S0 (nx36231)) ;
    mux21_ni ix15704 (.Y (nx15703), .A0 (label_3_output[9]), .A1 (
             label_3_input_9), .S0 (nx36269)) ;
    mux21_ni ix3365 (.Y (nx3364), .A0 (nx3360), .A1 (
             label_3_input_state_machine_9), .S0 (nx35947)) ;
    mux21_ni ix15694 (.Y (nx15693), .A0 (label_3_input_state_machine_9), .A1 (
             mdr_data_out[41]), .S0 (nx36231)) ;
    mux21_ni ix15664 (.Y (nx15663), .A0 (label_3_output[7]), .A1 (
             label_3_input_7), .S0 (nx36269)) ;
    mux21_ni ix3301 (.Y (nx3300), .A0 (nx3296), .A1 (
             label_3_input_state_machine_7), .S0 (nx35947)) ;
    mux21_ni ix15654 (.Y (nx15653), .A0 (label_3_input_state_machine_7), .A1 (
             mdr_data_out[39]), .S0 (nx36233)) ;
    mux21_ni ix15624 (.Y (nx15623), .A0 (label_3_output[5]), .A1 (
             label_3_input_5), .S0 (nx36271)) ;
    mux21_ni ix3237 (.Y (nx3236), .A0 (nx3232), .A1 (
             label_3_input_state_machine_5), .S0 (nx35169)) ;
    mux21_ni ix15614 (.Y (nx15613), .A0 (label_3_input_state_machine_5), .A1 (
             mdr_data_out[37]), .S0 (nx36233)) ;
    mux21_ni ix15584 (.Y (nx15583), .A0 (label_3_output[3]), .A1 (
             label_3_input_3), .S0 (nx36271)) ;
    mux21_ni ix3173 (.Y (nx3172), .A0 (nx3168), .A1 (
             label_3_input_state_machine_3), .S0 (nx35169)) ;
    mux21_ni ix15574 (.Y (nx15573), .A0 (label_3_input_state_machine_3), .A1 (
             mdr_data_out[35]), .S0 (nx36233)) ;
    mux21_ni ix15544 (.Y (nx15543), .A0 (label_3_output[1]), .A1 (
             label_3_input_1), .S0 (nx36271)) ;
    mux21_ni ix3109 (.Y (nx3108), .A0 (nx3104), .A1 (
             label_3_input_state_machine_1), .S0 (nx35169)) ;
    mux21_ni ix15534 (.Y (nx15533), .A0 (label_3_input_state_machine_1), .A1 (
             mdr_data_out[33]), .S0 (nx36233)) ;
    xnor2 ix32765 (.Y (nx32764), .A0 (nx29051), .A1 (nx32774)) ;
    mux21_ni ix15564 (.Y (nx15563), .A0 (label_3_output[2]), .A1 (
             label_3_input_2), .S0 (nx36271)) ;
    mux21_ni ix3141 (.Y (nx3140), .A0 (nx3136), .A1 (
             label_3_input_state_machine_2), .S0 (nx35169)) ;
    mux21_ni ix15554 (.Y (nx15553), .A0 (label_3_input_state_machine_2), .A1 (
             mdr_data_out[34]), .S0 (nx36233)) ;
    xnor2 ix32780 (.Y (nx32779), .A0 (nx29049), .A1 (nx32789)) ;
    mux21_ni ix15604 (.Y (nx15603), .A0 (label_3_output[4]), .A1 (
             label_3_input_4), .S0 (nx36271)) ;
    mux21_ni ix3205 (.Y (nx3204), .A0 (nx3200), .A1 (
             label_3_input_state_machine_4), .S0 (nx35169)) ;
    mux21_ni ix15594 (.Y (nx15593), .A0 (label_3_input_state_machine_4), .A1 (
             mdr_data_out[36]), .S0 (nx36233)) ;
    xnor2 ix32795 (.Y (nx32794), .A0 (nx29047), .A1 (nx32804)) ;
    mux21_ni ix15644 (.Y (nx15643), .A0 (label_3_output[6]), .A1 (
             label_3_input_6), .S0 (nx36271)) ;
    mux21_ni ix3269 (.Y (nx3268), .A0 (nx3264), .A1 (
             label_3_input_state_machine_6), .S0 (nx35169)) ;
    mux21_ni ix15634 (.Y (nx15633), .A0 (label_3_input_state_machine_6), .A1 (
             mdr_data_out[38]), .S0 (nx36233)) ;
    xnor2 ix32810 (.Y (nx32809), .A0 (nx29045), .A1 (nx32819)) ;
    mux21_ni ix15684 (.Y (nx15683), .A0 (label_3_output[8]), .A1 (
             label_3_input_8), .S0 (nx36271)) ;
    mux21_ni ix3333 (.Y (nx3332), .A0 (nx3328), .A1 (
             label_3_input_state_machine_8), .S0 (nx35169)) ;
    mux21_ni ix15674 (.Y (nx15673), .A0 (label_3_input_state_machine_8), .A1 (
             mdr_data_out[40]), .S0 (nx36235)) ;
    xnor2 ix32825 (.Y (nx32824), .A0 (nx29043), .A1 (nx32834)) ;
    mux21_ni ix15724 (.Y (nx15723), .A0 (label_3_output[10]), .A1 (
             label_3_input_10), .S0 (nx36273)) ;
    mux21_ni ix3397 (.Y (nx3396), .A0 (nx3392), .A1 (
             label_3_input_state_machine_10), .S0 (nx35949)) ;
    mux21_ni ix15714 (.Y (nx15713), .A0 (label_3_input_state_machine_10), .A1 (
             mdr_data_out[42]), .S0 (nx36235)) ;
    xnor2 ix32840 (.Y (nx32839), .A0 (nx29041), .A1 (nx32849)) ;
    mux21_ni ix15764 (.Y (nx15763), .A0 (label_3_output[12]), .A1 (
             label_3_input_12), .S0 (nx36273)) ;
    mux21_ni ix3461 (.Y (nx3460), .A0 (nx3456), .A1 (
             label_3_input_state_machine_12), .S0 (nx35949)) ;
    mux21_ni ix15754 (.Y (nx15753), .A0 (label_3_input_state_machine_12), .A1 (
             mdr_data_out[44]), .S0 (nx36235)) ;
    xnor2 ix32855 (.Y (nx32854), .A0 (nx29039), .A1 (nx32856)) ;
    ao32 ix21664 (.Y (nx21663), .A0 (nx35961), .A1 (nx35653), .A2 (nx36293), .B0 (
         max_calc_ans3_14), .B1 (nx35877)) ;
    mux21 ix32860 (.Y (nx35653), .A0 (nx29942), .A1 (nx30132), .S0 (nx35887)) ;
    xnor2 ix15909 (.Y (nx15908), .A0 (nx32472), .A1 (nx32669)) ;
    xnor2 ix32866 (.Y (nx32865), .A0 (nx32869), .A1 (
          max_calc_comparator_second_inp1_13)) ;
    mux21_ni ix15935 (.Y (nx15934), .A0 (max_calc_ans4_13), .A1 (
             label_4_output[13]), .S0 (nx35979)) ;
    ao32 ix23724 (.Y (nx23723), .A0 (nx35961), .A1 (nx35655), .A2 (nx36293), .B0 (
         max_calc_ans4_13), .B1 (nx35877)) ;
    mux21 ix32877 (.Y (nx35655), .A0 (nx32252), .A1 (nx32256), .S0 (nx35893)) ;
    mux21_ni ix15971 (.Y (nx15970), .A0 (max_calc_ans3_13), .A1 (
             label_3_output[13]), .S0 (nx35979)) ;
    ao32 ix23744 (.Y (nx23743), .A0 (nx35961), .A1 (nx35657), .A2 (nx36293), .B0 (
         max_calc_ans3_13), .B1 (nx35877)) ;
    mux21 ix32889 (.Y (nx35657), .A0 (nx30325), .A1 (nx30329), .S0 (nx35887)) ;
    mux21 ix16009 (.Y (nx16008), .A0 (nx32904), .A1 (nx32653), .S0 (nx35979)) ;
    ao32 ix23764 (.Y (nx23763), .A0 (nx35961), .A1 (nx35659), .A2 (nx36293), .B0 (
         max_calc_ans4_12), .B1 (nx35877)) ;
    mux21 ix32903 (.Y (nx35659), .A0 (nx32263), .A1 (nx32270), .S0 (nx35893)) ;
    mux21 ix16045 (.Y (nx16044), .A0 (nx32917), .A1 (nx32849), .S0 (nx35981)) ;
    ao32 ix23784 (.Y (nx23783), .A0 (nx35961), .A1 (nx35661), .A2 (nx36293), .B0 (
         max_calc_ans3_12), .B1 (nx35879)) ;
    mux21 ix32916 (.Y (nx35661), .A0 (nx30336), .A1 (nx30343), .S0 (nx35887)) ;
    xnor2 ix16057 (.Y (nx16056), .A0 (nx32894), .A1 (nx32908)) ;
    xnor2 ix32922 (.Y (nx32921), .A0 (nx32925), .A1 (
          max_calc_comparator_second_inp1_11)) ;
    mux21_ni ix16083 (.Y (nx16082), .A0 (max_calc_ans4_11), .A1 (
             label_4_output[11]), .S0 (nx35981)) ;
    ao32 ix23804 (.Y (nx23803), .A0 (nx35963), .A1 (nx35663), .A2 (nx36293), .B0 (
         max_calc_ans4_11), .B1 (nx35879)) ;
    mux21 ix32933 (.Y (nx35663), .A0 (nx32280), .A1 (nx32284), .S0 (nx35893)) ;
    mux21_ni ix16119 (.Y (nx16118), .A0 (max_calc_ans3_11), .A1 (
             label_3_output[11]), .S0 (nx35981)) ;
    ao32 ix23824 (.Y (nx23823), .A0 (nx35963), .A1 (nx35665), .A2 (nx36293), .B0 (
         max_calc_ans3_11), .B1 (nx35879)) ;
    mux21 ix32945 (.Y (nx35665), .A0 (nx30353), .A1 (nx30357), .S0 (nx35887)) ;
    mux21 ix16157 (.Y (nx16156), .A0 (nx32960), .A1 (nx32638), .S0 (nx35981)) ;
    ao32 ix23844 (.Y (nx23843), .A0 (nx35963), .A1 (nx35667), .A2 (nx36295), .B0 (
         max_calc_ans4_10), .B1 (nx35879)) ;
    mux21 ix32959 (.Y (nx35667), .A0 (nx32291), .A1 (nx32298), .S0 (nx35893)) ;
    mux21 ix16193 (.Y (nx16192), .A0 (nx32973), .A1 (nx32834), .S0 (nx35981)) ;
    ao32 ix23864 (.Y (nx23863), .A0 (nx35963), .A1 (nx35669), .A2 (nx36295), .B0 (
         max_calc_ans3_10), .B1 (nx35879)) ;
    mux21 ix32972 (.Y (nx35669), .A0 (nx30364), .A1 (nx30371), .S0 (nx35887)) ;
    xnor2 ix16205 (.Y (nx16204), .A0 (nx32950), .A1 (nx32964)) ;
    xnor2 ix32978 (.Y (nx32977), .A0 (nx32981), .A1 (
          max_calc_comparator_second_inp1_9)) ;
    mux21_ni ix16231 (.Y (nx16230), .A0 (max_calc_ans4_9), .A1 (
             label_4_output[9]), .S0 (nx35981)) ;
    ao32 ix23884 (.Y (nx23883), .A0 (nx35963), .A1 (nx35671), .A2 (nx36295), .B0 (
         max_calc_ans4_9), .B1 (nx35879)) ;
    mux21 ix32989 (.Y (nx35671), .A0 (nx32308), .A1 (nx32312), .S0 (nx35893)) ;
    mux21_ni ix16267 (.Y (nx16266), .A0 (max_calc_ans3_9), .A1 (
             label_3_output[9]), .S0 (nx35981)) ;
    ao32 ix23904 (.Y (nx23903), .A0 (nx35963), .A1 (nx35673), .A2 (nx36295), .B0 (
         max_calc_ans3_9), .B1 (nx35879)) ;
    mux21 ix33001 (.Y (nx35673), .A0 (nx30381), .A1 (nx30385), .S0 (nx35887)) ;
    mux21 ix16305 (.Y (nx16304), .A0 (nx33016), .A1 (nx32623), .S0 (nx35983)) ;
    ao32 ix23924 (.Y (nx23923), .A0 (nx35963), .A1 (nx35675), .A2 (nx36295), .B0 (
         max_calc_ans4_8), .B1 (nx35881)) ;
    mux21 ix33015 (.Y (nx35675), .A0 (nx32319), .A1 (nx32326), .S0 (nx35895)) ;
    mux21 ix16341 (.Y (nx16340), .A0 (nx33029), .A1 (nx32819), .S0 (nx35983)) ;
    ao32 ix23944 (.Y (nx23943), .A0 (nx35183), .A1 (nx35677), .A2 (nx36295), .B0 (
         max_calc_ans3_8), .B1 (nx35881)) ;
    mux21 ix33028 (.Y (nx35677), .A0 (nx30392), .A1 (nx30399), .S0 (nx35889)) ;
    xnor2 ix16353 (.Y (nx16352), .A0 (nx33006), .A1 (nx33020)) ;
    xnor2 ix33034 (.Y (nx33033), .A0 (nx33037), .A1 (
          max_calc_comparator_second_inp1_7)) ;
    mux21_ni ix16379 (.Y (nx16378), .A0 (max_calc_ans4_7), .A1 (
             label_4_output[7]), .S0 (nx35983)) ;
    ao32 ix23964 (.Y (nx23963), .A0 (nx35183), .A1 (nx35679), .A2 (nx36295), .B0 (
         max_calc_ans4_7), .B1 (nx35881)) ;
    mux21 ix33045 (.Y (nx35679), .A0 (nx32336), .A1 (nx32340), .S0 (nx35895)) ;
    mux21_ni ix16415 (.Y (nx16414), .A0 (max_calc_ans3_7), .A1 (
             label_3_output[7]), .S0 (nx35983)) ;
    ao32 ix23984 (.Y (nx23983), .A0 (nx35183), .A1 (nx35681), .A2 (nx36297), .B0 (
         max_calc_ans3_7), .B1 (nx35881)) ;
    mux21 ix33057 (.Y (nx35681), .A0 (nx30409), .A1 (nx30413), .S0 (nx35889)) ;
    mux21 ix16453 (.Y (nx16452), .A0 (nx33072), .A1 (nx32608), .S0 (nx35983)) ;
    ao32 ix24004 (.Y (nx24003), .A0 (nx35965), .A1 (nx35683), .A2 (nx36297), .B0 (
         max_calc_ans4_6), .B1 (nx35881)) ;
    mux21 ix33071 (.Y (nx35683), .A0 (nx32347), .A1 (nx32354), .S0 (nx35895)) ;
    mux21 ix16489 (.Y (nx16488), .A0 (nx33085), .A1 (nx32804), .S0 (nx35983)) ;
    ao32 ix24024 (.Y (nx24023), .A0 (nx35965), .A1 (nx35685), .A2 (nx36297), .B0 (
         max_calc_ans3_6), .B1 (nx35881)) ;
    mux21 ix33084 (.Y (nx35685), .A0 (nx30420), .A1 (nx30427), .S0 (nx35889)) ;
    xnor2 ix16501 (.Y (nx16500), .A0 (nx33062), .A1 (nx33076)) ;
    xnor2 ix33090 (.Y (nx33089), .A0 (nx33093), .A1 (
          max_calc_comparator_second_inp1_5)) ;
    mux21_ni ix16527 (.Y (nx16526), .A0 (max_calc_ans4_5), .A1 (
             label_4_output[5]), .S0 (nx35983)) ;
    ao32 ix24044 (.Y (nx24043), .A0 (nx35965), .A1 (nx35687), .A2 (nx36297), .B0 (
         max_calc_ans4_5), .B1 (nx35881)) ;
    mux21 ix33101 (.Y (nx35687), .A0 (nx32364), .A1 (nx32368), .S0 (nx35895)) ;
    mux21_ni ix16563 (.Y (nx16562), .A0 (max_calc_ans3_5), .A1 (
             label_3_output[5]), .S0 (nx35985)) ;
    ao32 ix24064 (.Y (nx24063), .A0 (nx35965), .A1 (nx35689), .A2 (nx36297), .B0 (
         max_calc_ans3_5), .B1 (nx35883)) ;
    mux21 ix33113 (.Y (nx35689), .A0 (nx30437), .A1 (nx30441), .S0 (nx35889)) ;
    mux21 ix16601 (.Y (nx16600), .A0 (nx33128), .A1 (nx32593), .S0 (nx35985)) ;
    ao32 ix24084 (.Y (nx24083), .A0 (nx35965), .A1 (nx35691), .A2 (nx36297), .B0 (
         max_calc_ans4_4), .B1 (nx35883)) ;
    mux21 ix33127 (.Y (nx35691), .A0 (nx32375), .A1 (nx32382), .S0 (nx35895)) ;
    mux21 ix16637 (.Y (nx16636), .A0 (nx33141), .A1 (nx32789), .S0 (nx35985)) ;
    ao32 ix24104 (.Y (nx24103), .A0 (nx35965), .A1 (nx35693), .A2 (nx36297), .B0 (
         max_calc_ans3_4), .B1 (nx35883)) ;
    mux21 ix33140 (.Y (nx35693), .A0 (nx30448), .A1 (nx30455), .S0 (nx35889)) ;
    xnor2 ix16649 (.Y (nx16648), .A0 (nx33118), .A1 (nx33132)) ;
    xnor2 ix33146 (.Y (nx33145), .A0 (nx33149), .A1 (
          max_calc_comparator_second_inp1_3)) ;
    mux21_ni ix16675 (.Y (nx16674), .A0 (max_calc_ans4_3), .A1 (
             label_4_output[3]), .S0 (nx35985)) ;
    ao32 ix24124 (.Y (nx24123), .A0 (nx35967), .A1 (nx35695), .A2 (nx36393), .B0 (
         max_calc_ans4_3), .B1 (nx35883)) ;
    mux21 ix33157 (.Y (nx35695), .A0 (nx32392), .A1 (nx32396), .S0 (nx35895)) ;
    mux21_ni ix16711 (.Y (nx16710), .A0 (max_calc_ans3_3), .A1 (
             label_3_output[3]), .S0 (nx35985)) ;
    ao32 ix24144 (.Y (nx24143), .A0 (nx35967), .A1 (nx35697), .A2 (nx36393), .B0 (
         max_calc_ans3_3), .B1 (nx35883)) ;
    mux21 ix33169 (.Y (nx35697), .A0 (nx30465), .A1 (nx30469), .S0 (nx35889)) ;
    mux21 ix16749 (.Y (nx16748), .A0 (nx33184), .A1 (nx32578), .S0 (nx35985)) ;
    ao32 ix24164 (.Y (nx24163), .A0 (nx35967), .A1 (nx35699), .A2 (nx36393), .B0 (
         max_calc_ans4_2), .B1 (nx35883)) ;
    mux21 ix33183 (.Y (nx35699), .A0 (nx32403), .A1 (nx32410), .S0 (nx35895)) ;
    mux21 ix16785 (.Y (nx16784), .A0 (nx33197), .A1 (nx32774), .S0 (nx35985)) ;
    ao32 ix24184 (.Y (nx24183), .A0 (nx35967), .A1 (nx35701), .A2 (nx36393), .B0 (
         max_calc_ans3_2), .B1 (nx35883)) ;
    mux21 ix33196 (.Y (nx35701), .A0 (nx30476), .A1 (nx30483), .S0 (nx35889)) ;
    xnor2 ix16797 (.Y (nx16796), .A0 (nx33174), .A1 (nx33188)) ;
    mux21_ni ix16823 (.Y (nx16822), .A0 (max_calc_ans4_1), .A1 (
             label_4_output[1]), .S0 (nx35187)) ;
    ao32 ix24204 (.Y (nx24203), .A0 (nx35967), .A1 (nx35703), .A2 (nx36393), .B0 (
         max_calc_ans4_1), .B1 (nx35885)) ;
    mux21 ix33211 (.Y (nx35703), .A0 (nx32418), .A1 (nx32422), .S0 (nx35897)) ;
    mux21_ni ix16859 (.Y (nx16858), .A0 (max_calc_ans3_1), .A1 (
             label_3_output[1]), .S0 (nx35987)) ;
    ao32 ix24224 (.Y (nx24223), .A0 (nx35967), .A1 (nx35705), .A2 (nx36393), .B0 (
         max_calc_ans3_1), .B1 (nx35885)) ;
    mux21 ix33223 (.Y (nx35705), .A0 (nx30491), .A1 (nx30495), .S0 (nx35891)) ;
    xnor2 ix16871 (.Y (nx16870), .A0 (nx33203), .A1 (nx33214)) ;
    xnor2 ix17137 (.Y (nx17136), .A0 (nx33232), .A1 (nx33257)) ;
    mux21_ni ix17089 (.Y (nx17088), .A0 (max_calc_ans4_15), .A1 (
             label_4_output[15]), .S0 (nx35987)) ;
    mux21_ni ix14964 (.Y (nx14963), .A0 (label_4_output[15]), .A1 (
             label_4_input_15), .S0 (nx36273)) ;
    mux21_ni ix2213 (.Y (nx2212), .A0 (nx2208), .A1 (
             label_4_input_state_machine_15), .S0 (nx35949)) ;
    mux21_ni ix14124 (.Y (nx14123), .A0 (label_4_input_state_machine_15), .A1 (
             mdr_data_out[63]), .S0 (nx36235)) ;
    xor2 ix33247 (.Y (nx33246), .A0 (nx30966), .A1 (label_4_output[15])) ;
    ao32 ix24284 (.Y (nx24283), .A0 (nx35967), .A1 (nx35707), .A2 (nx36393), .B0 (
         max_calc_ans4_15), .B1 (nx35885)) ;
    mux21 ix33252 (.Y (nx35707), .A0 (nx32433), .A1 (nx32451), .S0 (nx35897)) ;
    mux21_ni ix17125 (.Y (nx17124), .A0 (max_calc_ans3_15), .A1 (
             label_3_output[15]), .S0 (nx35987)) ;
    mux21_ni ix15814 (.Y (nx15813), .A0 (label_3_output[15]), .A1 (
             label_3_input_15), .S0 (nx36273)) ;
    mux21_ni ix3551 (.Y (nx3550), .A0 (nx3546), .A1 (
             label_3_input_state_machine_15), .S0 (nx35949)) ;
    mux21_ni ix14974 (.Y (nx14973), .A0 (label_3_input_state_machine_15), .A1 (
             mdr_data_out[47]), .S0 (nx36235)) ;
    xor2 ix33272 (.Y (nx33271), .A0 (nx29037), .A1 (label_3_output[15])) ;
    ao32 ix24304 (.Y (nx24303), .A0 (nx35969), .A1 (nx35709), .A2 (nx35749), .B0 (
         max_calc_ans3_15), .B1 (nx35885)) ;
    mux21 ix33277 (.Y (nx35709), .A0 (nx30506), .A1 (nx30524), .S0 (nx35891)) ;
    mux21_ni ix18889 (.Y (nx18888), .A0 (max_calc_ans8_0), .A1 (max_calc_ans7_0)
             , .S0 (nx35987)) ;
    mux21_ni ix25464 (.Y (nx25463), .A0 (max_calc_ans7_0), .A1 (nx18854), .S0 (
             nx36021)) ;
    mux21_ni ix25454 (.Y (nx25453), .A0 (nx13121), .A1 (max_calc_ans8_0), .S0 (
             nx35869)) ;
    mux21_ni ix24394 (.Y (nx24393), .A0 (max_calc_comparator_first_inp2_14), .A1 (
             nx17248), .S0 (nx36281)) ;
    mux21_ni ix17249 (.Y (nx17248), .A0 (nx17244), .A1 (nx17156), .S0 (nx35969)
             ) ;
    mux21_ni ix17157 (.Y (nx17156), .A0 (max_calc_ans2_14), .A1 (
             label_2_output[14]), .S0 (nx35987)) ;
    mux21_ni ix16654 (.Y (nx16653), .A0 (label_2_output[14]), .A1 (
             label_2_input_14), .S0 (nx36273)) ;
    mux21_ni ix4863 (.Y (nx4862), .A0 (nx4858), .A1 (
             label_2_input_state_machine_14), .S0 (nx35951)) ;
    mux21_ni ix16644 (.Y (nx16643), .A0 (label_2_input_state_machine_14), .A1 (
             mdr_data_out[30]), .S0 (nx36235)) ;
    mux21_ni ix16634 (.Y (nx16633), .A0 (label_2_output[13]), .A1 (
             label_2_input_13), .S0 (nx36273)) ;
    mux21_ni ix4831 (.Y (nx4830), .A0 (nx4826), .A1 (
             label_2_input_state_machine_13), .S0 (nx35951)) ;
    mux21_ni ix16624 (.Y (nx16623), .A0 (label_2_input_state_machine_13), .A1 (
             mdr_data_out[29]), .S0 (nx36235)) ;
    mux21_ni ix16594 (.Y (nx16593), .A0 (label_2_output[11]), .A1 (
             label_2_input_11), .S0 (nx36273)) ;
    mux21_ni ix4767 (.Y (nx4766), .A0 (nx4762), .A1 (
             label_2_input_state_machine_11), .S0 (nx35951)) ;
    mux21_ni ix16584 (.Y (nx16583), .A0 (label_2_input_state_machine_11), .A1 (
             mdr_data_out[27]), .S0 (nx35599)) ;
    mux21_ni ix16554 (.Y (nx16553), .A0 (label_2_output[9]), .A1 (
             label_2_input_9), .S0 (nx36275)) ;
    mux21_ni ix4703 (.Y (nx4702), .A0 (nx4698), .A1 (
             label_2_input_state_machine_9), .S0 (nx35951)) ;
    mux21_ni ix16544 (.Y (nx16543), .A0 (label_2_input_state_machine_9), .A1 (
             mdr_data_out[25]), .S0 (nx35599)) ;
    mux21_ni ix16514 (.Y (nx16513), .A0 (label_2_output[7]), .A1 (
             label_2_input_7), .S0 (nx36275)) ;
    mux21_ni ix4639 (.Y (nx4638), .A0 (nx4634), .A1 (
             label_2_input_state_machine_7), .S0 (nx35951)) ;
    mux21_ni ix16504 (.Y (nx16503), .A0 (label_2_input_state_machine_7), .A1 (
             mdr_data_out[23]), .S0 (nx35599)) ;
    mux21_ni ix16474 (.Y (nx16473), .A0 (label_2_output[5]), .A1 (
             label_2_input_5), .S0 (nx36275)) ;
    mux21_ni ix4575 (.Y (nx4574), .A0 (nx4570), .A1 (
             label_2_input_state_machine_5), .S0 (nx35951)) ;
    mux21_ni ix16464 (.Y (nx16463), .A0 (label_2_input_state_machine_5), .A1 (
             mdr_data_out[21]), .S0 (nx35599)) ;
    mux21_ni ix16434 (.Y (nx16433), .A0 (label_2_output[3]), .A1 (
             label_2_input_3), .S0 (nx36275)) ;
    mux21_ni ix4511 (.Y (nx4510), .A0 (nx4506), .A1 (
             label_2_input_state_machine_3), .S0 (nx35951)) ;
    mux21_ni ix16424 (.Y (nx16423), .A0 (label_2_input_state_machine_3), .A1 (
             mdr_data_out[19]), .S0 (nx35599)) ;
    mux21_ni ix16394 (.Y (nx16393), .A0 (label_2_output[1]), .A1 (
             label_2_input_1), .S0 (nx36275)) ;
    mux21_ni ix4447 (.Y (nx4446), .A0 (nx4442), .A1 (
             label_2_input_state_machine_1), .S0 (nx35953)) ;
    mux21_ni ix16384 (.Y (nx16383), .A0 (label_2_input_state_machine_1), .A1 (
             mdr_data_out[17]), .S0 (nx35599)) ;
    xnor2 ix33388 (.Y (nx33387), .A0 (nx28608), .A1 (nx33397)) ;
    mux21_ni ix16414 (.Y (nx16413), .A0 (label_2_output[2]), .A1 (
             label_2_input_2), .S0 (nx36275)) ;
    mux21_ni ix4479 (.Y (nx4478), .A0 (nx4474), .A1 (
             label_2_input_state_machine_2), .S0 (nx35953)) ;
    mux21_ni ix16404 (.Y (nx16403), .A0 (label_2_input_state_machine_2), .A1 (
             mdr_data_out[18]), .S0 (nx35599)) ;
    xnor2 ix33403 (.Y (nx33402), .A0 (nx28606), .A1 (nx33412)) ;
    mux21_ni ix16454 (.Y (nx16453), .A0 (label_2_output[4]), .A1 (
             label_2_input_4), .S0 (nx36275)) ;
    mux21_ni ix4543 (.Y (nx4542), .A0 (nx4538), .A1 (
             label_2_input_state_machine_4), .S0 (nx35953)) ;
    mux21_ni ix16444 (.Y (nx16443), .A0 (label_2_input_state_machine_4), .A1 (
             mdr_data_out[20]), .S0 (nx36237)) ;
    xnor2 ix33418 (.Y (nx33417), .A0 (nx28604), .A1 (nx33427)) ;
    mux21_ni ix16494 (.Y (nx16493), .A0 (label_2_output[6]), .A1 (
             label_2_input_6), .S0 (nx35607)) ;
    mux21_ni ix4607 (.Y (nx4606), .A0 (nx4602), .A1 (
             label_2_input_state_machine_6), .S0 (nx35953)) ;
    mux21_ni ix16484 (.Y (nx16483), .A0 (label_2_input_state_machine_6), .A1 (
             mdr_data_out[22]), .S0 (nx36237)) ;
    xnor2 ix33433 (.Y (nx33432), .A0 (nx28602), .A1 (nx33442)) ;
    mux21_ni ix16534 (.Y (nx16533), .A0 (label_2_output[8]), .A1 (
             label_2_input_8), .S0 (nx35607)) ;
    mux21_ni ix4671 (.Y (nx4670), .A0 (nx4666), .A1 (
             label_2_input_state_machine_8), .S0 (nx35953)) ;
    mux21_ni ix16524 (.Y (nx16523), .A0 (label_2_input_state_machine_8), .A1 (
             mdr_data_out[24]), .S0 (nx36237)) ;
    xnor2 ix33448 (.Y (nx33447), .A0 (nx28600), .A1 (nx33457)) ;
    mux21_ni ix16574 (.Y (nx16573), .A0 (label_2_output[10]), .A1 (
             label_2_input_10), .S0 (nx35607)) ;
    mux21_ni ix4735 (.Y (nx4734), .A0 (nx4730), .A1 (
             label_2_input_state_machine_10), .S0 (nx35953)) ;
    mux21_ni ix16564 (.Y (nx16563), .A0 (label_2_input_state_machine_10), .A1 (
             mdr_data_out[26]), .S0 (nx36237)) ;
    xnor2 ix33463 (.Y (nx33462), .A0 (nx28598), .A1 (nx33472)) ;
    mux21_ni ix16614 (.Y (nx16613), .A0 (label_2_output[12]), .A1 (
             label_2_input_12), .S0 (nx35607)) ;
    mux21_ni ix4799 (.Y (nx4798), .A0 (nx4794), .A1 (
             label_2_input_state_machine_12), .S0 (nx35953)) ;
    mux21_ni ix16604 (.Y (nx16603), .A0 (label_2_input_state_machine_12), .A1 (
             mdr_data_out[28]), .S0 (nx36237)) ;
    xnor2 ix33478 (.Y (nx33477), .A0 (nx28596), .A1 (nx33479)) ;
    mux21_ni ix24324 (.Y (nx24323), .A0 (nx17146), .A1 (max_calc_ans2_14), .S0 (
             nx35851)) ;
    mux21 ix17147 (.Y (nx17146), .A0 (nx32472), .A1 (nx32669), .S0 (nx35899)) ;
    mux21_ni ix17245 (.Y (nx17244), .A0 (max_calc_ans8_14), .A1 (
             max_calc_ans7_14), .S0 (nx35987)) ;
    mux21_ni ix24384 (.Y (nx24383), .A0 (max_calc_ans7_14), .A1 (nx17146), .S0 (
             nx36021)) ;
    mux21_ni ix24374 (.Y (nx24373), .A0 (nx13371), .A1 (max_calc_ans8_14), .S0 (
             nx35869)) ;
    mux21_ni ix17225 (.Y (nx13371), .A0 (max_calc_comparator_first_inp2_14), .A1 (
             max_calc_comparator_first_inp1_14), .S0 (nx35905)) ;
    mux21_ni ix24364 (.Y (nx24363), .A0 (max_calc_comparator_first_inp1_14), .A1 (
             nx17210), .S0 (nx36281)) ;
    mux21_ni ix17211 (.Y (nx17210), .A0 (nx17206), .A1 (nx17174), .S0 (nx35969)
             ) ;
    mux21_ni ix17175 (.Y (nx17174), .A0 (max_calc_ans1_14), .A1 (
             label_1_output[14]), .S0 (nx35989)) ;
    mux21_ni ix17504 (.Y (nx17503), .A0 (label_1_output[14]), .A1 (
             label_1_input_14), .S0 (nx36277)) ;
    mux21_ni ix6201 (.Y (nx6200), .A0 (nx6196), .A1 (
             label_1_input_state_machine_14), .S0 (nx35955)) ;
    mux21_ni ix17494 (.Y (nx17493), .A0 (label_1_input_state_machine_14), .A1 (
             mdr_data_out[14]), .S0 (nx36237)) ;
    mux21_ni ix17484 (.Y (nx17483), .A0 (label_1_output[13]), .A1 (
             label_1_input_13), .S0 (nx36277)) ;
    mux21_ni ix6169 (.Y (nx6168), .A0 (nx6164), .A1 (
             label_1_input_state_machine_13), .S0 (nx35955)) ;
    mux21_ni ix17474 (.Y (nx17473), .A0 (label_1_input_state_machine_13), .A1 (
             mdr_data_out[13]), .S0 (nx36237)) ;
    mux21_ni ix17444 (.Y (nx17443), .A0 (label_1_output[11]), .A1 (
             label_1_input_11), .S0 (nx36279)) ;
    mux21_ni ix6105 (.Y (nx6104), .A0 (nx6100), .A1 (
             label_1_input_state_machine_11), .S0 (nx35955)) ;
    mux21_ni ix17434 (.Y (nx17433), .A0 (label_1_input_state_machine_11), .A1 (
             mdr_data_out[11]), .S0 (nx36239)) ;
    mux21_ni ix17404 (.Y (nx17403), .A0 (label_1_output[9]), .A1 (
             label_1_input_9), .S0 (nx36279)) ;
    mux21_ni ix6041 (.Y (nx6040), .A0 (nx6036), .A1 (
             label_1_input_state_machine_9), .S0 (nx35955)) ;
    mux21_ni ix17394 (.Y (nx17393), .A0 (label_1_input_state_machine_9), .A1 (
             mdr_data_out[9]), .S0 (nx36239)) ;
    mux21_ni ix17364 (.Y (nx17363), .A0 (label_1_output[7]), .A1 (
             label_1_input_7), .S0 (nx36279)) ;
    mux21_ni ix5977 (.Y (nx5976), .A0 (nx5972), .A1 (
             label_1_input_state_machine_7), .S0 (nx35955)) ;
    mux21_ni ix17354 (.Y (nx17353), .A0 (label_1_input_state_machine_7), .A1 (
             mdr_data_out[7]), .S0 (nx36239)) ;
    mux21_ni ix17324 (.Y (nx17323), .A0 (label_1_output[5]), .A1 (
             label_1_input_5), .S0 (nx36279)) ;
    mux21_ni ix5913 (.Y (nx5912), .A0 (nx5908), .A1 (
             label_1_input_state_machine_5), .S0 (nx35955)) ;
    mux21_ni ix17314 (.Y (nx17313), .A0 (label_1_input_state_machine_5), .A1 (
             mdr_data_out[5]), .S0 (nx36239)) ;
    mux21_ni ix17284 (.Y (nx17283), .A0 (label_1_output[3]), .A1 (
             label_1_input_3), .S0 (nx35607)) ;
    mux21_ni ix5849 (.Y (nx5848), .A0 (nx5844), .A1 (
             label_1_input_state_machine_3), .S0 (nx35955)) ;
    mux21_ni ix17274 (.Y (nx17273), .A0 (label_1_input_state_machine_3), .A1 (
             mdr_data_out[3]), .S0 (nx36239)) ;
    mux21_ni ix17244 (.Y (nx17243), .A0 (label_1_output[1]), .A1 (
             label_1_input_1), .S0 (nx35607)) ;
    mux21_ni ix5785 (.Y (nx5784), .A0 (nx5780), .A1 (
             label_1_input_state_machine_1), .S0 (nx35957)) ;
    mux21_ni ix17234 (.Y (nx17233), .A0 (label_1_input_state_machine_1), .A1 (
             mdr_data_out[1]), .S0 (nx36239)) ;
    xnor2 ix33586 (.Y (nx33585), .A0 (nx26648), .A1 (nx33595)) ;
    mux21_ni ix17264 (.Y (nx17263), .A0 (label_1_output[2]), .A1 (
             label_1_input_2), .S0 (nx35607)) ;
    mux21_ni ix5817 (.Y (nx5816), .A0 (nx5812), .A1 (
             label_1_input_state_machine_2), .S0 (nx35957)) ;
    mux21_ni ix17254 (.Y (nx17253), .A0 (label_1_input_state_machine_2), .A1 (
             mdr_data_out[2]), .S0 (nx36239)) ;
    xnor2 ix33601 (.Y (nx33600), .A0 (nx26646), .A1 (nx33610)) ;
    mux21_ni ix17304 (.Y (nx17303), .A0 (label_1_output[4]), .A1 (
             label_1_input_4), .S0 (nx36279)) ;
    mux21_ni ix5881 (.Y (nx5880), .A0 (nx5876), .A1 (
             label_1_input_state_machine_4), .S0 (nx35957)) ;
    mux21_ni ix17294 (.Y (nx17293), .A0 (label_1_input_state_machine_4), .A1 (
             mdr_data_out[4]), .S0 (nx35601)) ;
    xnor2 ix33616 (.Y (nx33615), .A0 (nx26644), .A1 (nx33625)) ;
    mux21_ni ix17344 (.Y (nx17343), .A0 (label_1_output[6]), .A1 (
             label_1_input_6), .S0 (nx36279)) ;
    mux21_ni ix5945 (.Y (nx5944), .A0 (nx5940), .A1 (
             label_1_input_state_machine_6), .S0 (nx35957)) ;
    mux21_ni ix17334 (.Y (nx17333), .A0 (label_1_input_state_machine_6), .A1 (
             mdr_data_out[6]), .S0 (nx35601)) ;
    xnor2 ix33631 (.Y (nx33630), .A0 (nx26642), .A1 (nx33640)) ;
    mux21_ni ix17384 (.Y (nx17383), .A0 (label_1_output[8]), .A1 (
             label_1_input_8), .S0 (nx36279)) ;
    mux21_ni ix6009 (.Y (nx6008), .A0 (nx6004), .A1 (
             label_1_input_state_machine_8), .S0 (nx35957)) ;
    mux21_ni ix17374 (.Y (nx17373), .A0 (label_1_input_state_machine_8), .A1 (
             mdr_data_out[8]), .S0 (nx35601)) ;
    xnor2 ix33646 (.Y (nx33645), .A0 (nx26640), .A1 (nx33655)) ;
    mux21_ni ix17424 (.Y (nx17423), .A0 (label_1_output[10]), .A1 (
             label_1_input_10), .S0 (nx35609)) ;
    mux21_ni ix6073 (.Y (nx6072), .A0 (nx6068), .A1 (
             label_1_input_state_machine_10), .S0 (nx35957)) ;
    mux21_ni ix17414 (.Y (nx17413), .A0 (label_1_input_state_machine_10), .A1 (
             mdr_data_out[10]), .S0 (nx35601)) ;
    xnor2 ix33661 (.Y (nx33660), .A0 (nx26638), .A1 (nx33670)) ;
    mux21_ni ix17464 (.Y (nx17463), .A0 (label_1_output[12]), .A1 (
             label_1_input_12), .S0 (nx35609)) ;
    mux21_ni ix6137 (.Y (nx6136), .A0 (nx6132), .A1 (
             label_1_input_state_machine_12), .S0 (nx35957)) ;
    mux21_ni ix17454 (.Y (nx17453), .A0 (label_1_input_state_machine_12), .A1 (
             mdr_data_out[12]), .S0 (nx35601)) ;
    xnor2 ix33676 (.Y (nx33675), .A0 (nx26636), .A1 (nx33677)) ;
    mux21_ni ix24334 (.Y (nx24333), .A0 (nx13371), .A1 (max_calc_ans1_14), .S0 (
             nx35851)) ;
    mux21_ni ix17207 (.Y (nx17206), .A0 (max_calc_ans5_14), .A1 (
             max_calc_ans6_14), .S0 (nx35989)) ;
    mux21_ni ix24344 (.Y (nx24343), .A0 (max_calc_ans6_14), .A1 (nx13371), .S0 (
             nx36021)) ;
    mux21_ni ix24354 (.Y (nx24353), .A0 (max_calc_ans5_14), .A1 (nx17196), .S0 (
             nx35749)) ;
    mux21 ix17197 (.Y (nx17196), .A0 (nx27573), .A1 (nx27763), .S0 (nx35861)) ;
    xor2 ix17257 (.Y (nx17256), .A0 (nx33292), .A1 (
         max_calc_comparator_first_inp1_14)) ;
    xor2 ix33695 (.Y (nx33694), .A0 (max_calc_comparator_first_inp2_13), .A1 (
         max_calc_comparator_first_inp1_13)) ;
    mux21_ni ix24474 (.Y (nx24473), .A0 (max_calc_comparator_first_inp2_13), .A1 (
             nx17370), .S0 (nx36281)) ;
    mux21_ni ix17371 (.Y (nx17370), .A0 (nx17366), .A1 (nx17278), .S0 (nx35969)
             ) ;
    mux21_ni ix17279 (.Y (nx17278), .A0 (max_calc_ans2_13), .A1 (
             label_2_output[13]), .S0 (nx35989)) ;
    mux21_ni ix24404 (.Y (nx24403), .A0 (nx17268), .A1 (max_calc_ans2_13), .S0 (
             nx35851)) ;
    mux21 ix17269 (.Y (nx17268), .A0 (nx32869), .A1 (nx32880), .S0 (nx35899)) ;
    mux21_ni ix17367 (.Y (nx17366), .A0 (max_calc_ans8_13), .A1 (
             max_calc_ans7_13), .S0 (nx35989)) ;
    mux21_ni ix24464 (.Y (nx24463), .A0 (max_calc_ans7_13), .A1 (nx17268), .S0 (
             nx36021)) ;
    mux21_ni ix24454 (.Y (nx24453), .A0 (nx13375), .A1 (max_calc_ans8_13), .S0 (
             nx35869)) ;
    mux21_ni ix17347 (.Y (nx13375), .A0 (max_calc_comparator_first_inp2_13), .A1 (
             max_calc_comparator_first_inp1_13), .S0 (nx35905)) ;
    mux21_ni ix24444 (.Y (nx24443), .A0 (max_calc_comparator_first_inp1_13), .A1 (
             nx17332), .S0 (nx36281)) ;
    mux21_ni ix17333 (.Y (nx17332), .A0 (nx17328), .A1 (nx17296), .S0 (nx35969)
             ) ;
    mux21_ni ix17297 (.Y (nx17296), .A0 (max_calc_ans1_13), .A1 (
             label_1_output[13]), .S0 (nx35989)) ;
    mux21_ni ix24414 (.Y (nx24413), .A0 (nx13375), .A1 (max_calc_ans1_13), .S0 (
             nx35851)) ;
    mux21_ni ix17329 (.Y (nx17328), .A0 (max_calc_ans5_13), .A1 (
             max_calc_ans6_13), .S0 (nx35989)) ;
    mux21_ni ix24424 (.Y (nx24423), .A0 (max_calc_ans6_13), .A1 (nx13375), .S0 (
             nx36021)) ;
    mux21_ni ix24434 (.Y (nx24433), .A0 (max_calc_ans5_13), .A1 (nx17318), .S0 (
             nx35749)) ;
    mux21 ix17319 (.Y (nx17318), .A0 (nx27956), .A1 (nx27960), .S0 (nx35861)) ;
    mux21_ni ix24554 (.Y (nx24553), .A0 (max_calc_comparator_first_inp2_12), .A1 (
             nx17492), .S0 (nx36283)) ;
    mux21_ni ix17493 (.Y (nx17492), .A0 (nx17488), .A1 (nx17400), .S0 (nx35969)
             ) ;
    mux21_ni ix17401 (.Y (nx17400), .A0 (max_calc_ans2_12), .A1 (
             label_2_output[12]), .S0 (nx35989)) ;
    mux21_ni ix24484 (.Y (nx24483), .A0 (nx17390), .A1 (max_calc_ans2_12), .S0 (
             nx35851)) ;
    mux21 ix17391 (.Y (nx17390), .A0 (nx32894), .A1 (nx32908), .S0 (nx35899)) ;
    mux21_ni ix17489 (.Y (nx17488), .A0 (max_calc_ans8_12), .A1 (
             max_calc_ans7_12), .S0 (nx35991)) ;
    mux21_ni ix24544 (.Y (nx24543), .A0 (max_calc_ans7_12), .A1 (nx17390), .S0 (
             nx36021)) ;
    mux21_ni ix24534 (.Y (nx24533), .A0 (nx13376), .A1 (max_calc_ans8_12), .S0 (
             nx35869)) ;
    mux21_ni ix17469 (.Y (nx13376), .A0 (max_calc_comparator_first_inp2_12), .A1 (
             max_calc_comparator_first_inp1_12), .S0 (nx35905)) ;
    mux21_ni ix24524 (.Y (nx24523), .A0 (max_calc_comparator_first_inp1_12), .A1 (
             nx17454), .S0 (nx36283)) ;
    mux21_ni ix17455 (.Y (nx17454), .A0 (nx17450), .A1 (nx17418), .S0 (nx35969)
             ) ;
    mux21_ni ix17419 (.Y (nx17418), .A0 (max_calc_ans1_12), .A1 (
             label_1_output[12]), .S0 (nx35991)) ;
    mux21_ni ix24494 (.Y (nx24493), .A0 (nx13376), .A1 (max_calc_ans1_12), .S0 (
             nx35853)) ;
    mux21_ni ix17451 (.Y (nx17450), .A0 (max_calc_ans5_12), .A1 (
             max_calc_ans6_12), .S0 (nx35991)) ;
    mux21_ni ix24504 (.Y (nx24503), .A0 (max_calc_ans6_12), .A1 (nx13376), .S0 (
             nx36023)) ;
    mux21_ni ix24514 (.Y (nx24513), .A0 (max_calc_ans5_12), .A1 (nx17440), .S0 (
             nx35749)) ;
    mux21 ix17441 (.Y (nx17440), .A0 (nx27967), .A1 (nx27974), .S0 (nx35861)) ;
    xor2 ix17501 (.Y (nx17500), .A0 (nx33731), .A1 (
         max_calc_comparator_first_inp1_12)) ;
    xor2 ix33768 (.Y (nx33767), .A0 (max_calc_comparator_first_inp2_11), .A1 (
         max_calc_comparator_first_inp1_11)) ;
    mux21_ni ix24634 (.Y (nx24633), .A0 (max_calc_comparator_first_inp2_11), .A1 (
             nx17614), .S0 (nx36283)) ;
    mux21_ni ix17615 (.Y (nx17614), .A0 (nx17610), .A1 (nx17522), .S0 (nx35971)
             ) ;
    mux21_ni ix17523 (.Y (nx17522), .A0 (max_calc_ans2_11), .A1 (
             label_2_output[11]), .S0 (nx35991)) ;
    mux21_ni ix24564 (.Y (nx24563), .A0 (nx17512), .A1 (max_calc_ans2_11), .S0 (
             nx35853)) ;
    mux21 ix17513 (.Y (nx17512), .A0 (nx32925), .A1 (nx32936), .S0 (nx35899)) ;
    mux21_ni ix17611 (.Y (nx17610), .A0 (max_calc_ans8_11), .A1 (
             max_calc_ans7_11), .S0 (nx35991)) ;
    mux21_ni ix24624 (.Y (nx24623), .A0 (max_calc_ans7_11), .A1 (nx17512), .S0 (
             nx36023)) ;
    mux21_ni ix24614 (.Y (nx24613), .A0 (nx13377), .A1 (max_calc_ans8_11), .S0 (
             nx35869)) ;
    mux21_ni ix17591 (.Y (nx13377), .A0 (max_calc_comparator_first_inp2_11), .A1 (
             max_calc_comparator_first_inp1_11), .S0 (nx35905)) ;
    mux21_ni ix24604 (.Y (nx24603), .A0 (max_calc_comparator_first_inp1_11), .A1 (
             nx17576), .S0 (nx36283)) ;
    mux21_ni ix17577 (.Y (nx17576), .A0 (nx17572), .A1 (nx17540), .S0 (nx35971)
             ) ;
    mux21_ni ix17541 (.Y (nx17540), .A0 (max_calc_ans1_11), .A1 (
             label_1_output[11]), .S0 (nx35991)) ;
    mux21_ni ix24574 (.Y (nx24573), .A0 (nx13377), .A1 (max_calc_ans1_11), .S0 (
             nx35853)) ;
    mux21_ni ix17573 (.Y (nx17572), .A0 (max_calc_ans5_11), .A1 (
             max_calc_ans6_11), .S0 (nx35991)) ;
    mux21_ni ix24584 (.Y (nx24583), .A0 (max_calc_ans6_11), .A1 (nx13377), .S0 (
             nx36023)) ;
    mux21_ni ix24594 (.Y (nx24593), .A0 (max_calc_ans5_11), .A1 (nx17562), .S0 (
             nx35749)) ;
    mux21 ix17563 (.Y (nx17562), .A0 (nx27984), .A1 (nx27988), .S0 (nx35861)) ;
    mux21_ni ix24714 (.Y (nx24713), .A0 (max_calc_comparator_first_inp2_10), .A1 (
             nx17736), .S0 (nx36283)) ;
    mux21_ni ix17737 (.Y (nx17736), .A0 (nx17732), .A1 (nx17644), .S0 (nx35971)
             ) ;
    mux21_ni ix17645 (.Y (nx17644), .A0 (max_calc_ans2_10), .A1 (
             label_2_output[10]), .S0 (nx35993)) ;
    mux21_ni ix24644 (.Y (nx24643), .A0 (nx17634), .A1 (max_calc_ans2_10), .S0 (
             nx35853)) ;
    mux21 ix17635 (.Y (nx17634), .A0 (nx32950), .A1 (nx32964), .S0 (nx35899)) ;
    mux21_ni ix17733 (.Y (nx17732), .A0 (max_calc_ans8_10), .A1 (
             max_calc_ans7_10), .S0 (nx35993)) ;
    mux21_ni ix24704 (.Y (nx24703), .A0 (max_calc_ans7_10), .A1 (nx17634), .S0 (
             nx36023)) ;
    mux21_ni ix24694 (.Y (nx24693), .A0 (nx13379), .A1 (max_calc_ans8_10), .S0 (
             nx35869)) ;
    mux21_ni ix17713 (.Y (nx13379), .A0 (max_calc_comparator_first_inp2_10), .A1 (
             max_calc_comparator_first_inp1_10), .S0 (nx35905)) ;
    mux21_ni ix24684 (.Y (nx24683), .A0 (max_calc_comparator_first_inp1_10), .A1 (
             nx17698), .S0 (nx36283)) ;
    mux21_ni ix17699 (.Y (nx17698), .A0 (nx17694), .A1 (nx17662), .S0 (nx35971)
             ) ;
    mux21_ni ix17663 (.Y (nx17662), .A0 (max_calc_ans1_10), .A1 (
             label_1_output[10]), .S0 (nx35993)) ;
    mux21_ni ix24654 (.Y (nx24653), .A0 (nx13379), .A1 (max_calc_ans1_10), .S0 (
             nx35853)) ;
    mux21_ni ix17695 (.Y (nx17694), .A0 (max_calc_ans5_10), .A1 (
             max_calc_ans6_10), .S0 (nx35993)) ;
    mux21_ni ix24664 (.Y (nx24663), .A0 (max_calc_ans6_10), .A1 (nx13379), .S0 (
             nx36023)) ;
    mux21_ni ix24674 (.Y (nx24673), .A0 (max_calc_ans5_10), .A1 (nx17684), .S0 (
             nx35749)) ;
    mux21 ix17685 (.Y (nx17684), .A0 (nx27995), .A1 (nx28002), .S0 (nx35861)) ;
    xor2 ix17745 (.Y (nx17744), .A0 (nx33804), .A1 (
         max_calc_comparator_first_inp1_10)) ;
    xor2 ix33841 (.Y (nx33840), .A0 (max_calc_comparator_first_inp2_9), .A1 (
         max_calc_comparator_first_inp1_9)) ;
    mux21_ni ix24794 (.Y (nx24793), .A0 (max_calc_comparator_first_inp2_9), .A1 (
             nx17858), .S0 (nx36283)) ;
    mux21_ni ix17859 (.Y (nx17858), .A0 (nx17854), .A1 (nx17766), .S0 (nx35971)
             ) ;
    mux21_ni ix17767 (.Y (nx17766), .A0 (max_calc_ans2_9), .A1 (
             label_2_output[9]), .S0 (nx35993)) ;
    mux21_ni ix24724 (.Y (nx24723), .A0 (nx17756), .A1 (max_calc_ans2_9), .S0 (
             nx35853)) ;
    mux21 ix17757 (.Y (nx17756), .A0 (nx32981), .A1 (nx32992), .S0 (nx35899)) ;
    mux21_ni ix17855 (.Y (nx17854), .A0 (max_calc_ans8_9), .A1 (max_calc_ans7_9)
             , .S0 (nx35993)) ;
    mux21_ni ix24784 (.Y (nx24783), .A0 (max_calc_ans7_9), .A1 (nx17756), .S0 (
             nx36023)) ;
    mux21_ni ix24774 (.Y (nx24773), .A0 (nx13381), .A1 (max_calc_ans8_9), .S0 (
             nx35871)) ;
    mux21_ni ix17835 (.Y (nx13381), .A0 (max_calc_comparator_first_inp2_9), .A1 (
             max_calc_comparator_first_inp1_9), .S0 (nx35905)) ;
    mux21_ni ix24764 (.Y (nx24763), .A0 (max_calc_comparator_first_inp1_9), .A1 (
             nx17820), .S0 (nx36285)) ;
    mux21_ni ix17821 (.Y (nx17820), .A0 (nx17816), .A1 (nx17784), .S0 (nx35971)
             ) ;
    mux21_ni ix17785 (.Y (nx17784), .A0 (max_calc_ans1_9), .A1 (
             label_1_output[9]), .S0 (nx35993)) ;
    mux21_ni ix24734 (.Y (nx24733), .A0 (nx13381), .A1 (max_calc_ans1_9), .S0 (
             nx35853)) ;
    mux21_ni ix17817 (.Y (nx17816), .A0 (max_calc_ans5_9), .A1 (max_calc_ans6_9)
             , .S0 (nx35995)) ;
    mux21_ni ix24744 (.Y (nx24743), .A0 (max_calc_ans6_9), .A1 (nx13381), .S0 (
             nx36023)) ;
    mux21_ni ix24754 (.Y (nx24753), .A0 (max_calc_ans5_9), .A1 (nx17806), .S0 (
             nx35749)) ;
    mux21 ix17807 (.Y (nx17806), .A0 (nx28012), .A1 (nx28016), .S0 (nx35861)) ;
    mux21_ni ix24874 (.Y (nx24873), .A0 (max_calc_comparator_first_inp2_8), .A1 (
             nx17980), .S0 (nx36285)) ;
    mux21_ni ix17981 (.Y (nx17980), .A0 (nx17976), .A1 (nx17888), .S0 (nx35971)
             ) ;
    mux21_ni ix17889 (.Y (nx17888), .A0 (max_calc_ans2_8), .A1 (
             label_2_output[8]), .S0 (nx35995)) ;
    mux21_ni ix24804 (.Y (nx24803), .A0 (nx17878), .A1 (max_calc_ans2_8), .S0 (
             nx35855)) ;
    mux21 ix17879 (.Y (nx17878), .A0 (nx33006), .A1 (nx33020), .S0 (nx35901)) ;
    mux21_ni ix17977 (.Y (nx17976), .A0 (max_calc_ans8_8), .A1 (max_calc_ans7_8)
             , .S0 (nx35995)) ;
    mux21_ni ix24864 (.Y (nx24863), .A0 (max_calc_ans7_8), .A1 (nx17878), .S0 (
             nx36025)) ;
    mux21_ni ix24854 (.Y (nx24853), .A0 (nx13383), .A1 (max_calc_ans8_8), .S0 (
             nx35871)) ;
    mux21_ni ix17957 (.Y (nx13383), .A0 (max_calc_comparator_first_inp2_8), .A1 (
             max_calc_comparator_first_inp1_8), .S0 (nx35907)) ;
    mux21_ni ix24844 (.Y (nx24843), .A0 (max_calc_comparator_first_inp1_8), .A1 (
             nx17942), .S0 (nx36285)) ;
    mux21_ni ix17943 (.Y (nx17942), .A0 (nx17938), .A1 (nx17906), .S0 (nx35973)
             ) ;
    mux21_ni ix17907 (.Y (nx17906), .A0 (max_calc_ans1_8), .A1 (
             label_1_output[8]), .S0 (nx35995)) ;
    mux21_ni ix24814 (.Y (nx24813), .A0 (nx13383), .A1 (max_calc_ans1_8), .S0 (
             nx35855)) ;
    mux21_ni ix17939 (.Y (nx17938), .A0 (max_calc_ans5_8), .A1 (max_calc_ans6_8)
             , .S0 (nx35995)) ;
    mux21_ni ix24824 (.Y (nx24823), .A0 (max_calc_ans6_8), .A1 (nx13383), .S0 (
             nx36025)) ;
    mux21_ni ix24834 (.Y (nx24833), .A0 (max_calc_ans5_8), .A1 (nx17928), .S0 (
             nx35751)) ;
    mux21 ix17929 (.Y (nx17928), .A0 (nx28023), .A1 (nx28030), .S0 (nx35863)) ;
    xor2 ix17989 (.Y (nx17988), .A0 (nx33877), .A1 (
         max_calc_comparator_first_inp1_8)) ;
    xor2 ix33914 (.Y (nx33913), .A0 (max_calc_comparator_first_inp2_7), .A1 (
         max_calc_comparator_first_inp1_7)) ;
    mux21_ni ix24954 (.Y (nx24953), .A0 (max_calc_comparator_first_inp2_7), .A1 (
             nx18102), .S0 (nx36285)) ;
    mux21_ni ix18103 (.Y (nx18102), .A0 (nx18098), .A1 (nx18010), .S0 (nx35973)
             ) ;
    mux21_ni ix18011 (.Y (nx18010), .A0 (max_calc_ans2_7), .A1 (
             label_2_output[7]), .S0 (nx35995)) ;
    mux21_ni ix24884 (.Y (nx24883), .A0 (nx18000), .A1 (max_calc_ans2_7), .S0 (
             nx35855)) ;
    mux21 ix18001 (.Y (nx18000), .A0 (nx33037), .A1 (nx33048), .S0 (nx35901)) ;
    mux21_ni ix18099 (.Y (nx18098), .A0 (max_calc_ans8_7), .A1 (max_calc_ans7_7)
             , .S0 (nx35995)) ;
    mux21_ni ix24944 (.Y (nx24943), .A0 (max_calc_ans7_7), .A1 (nx18000), .S0 (
             nx36025)) ;
    mux21_ni ix24934 (.Y (nx24933), .A0 (nx13385), .A1 (max_calc_ans8_7), .S0 (
             nx35871)) ;
    mux21_ni ix18079 (.Y (nx13385), .A0 (max_calc_comparator_first_inp2_7), .A1 (
             max_calc_comparator_first_inp1_7), .S0 (nx35907)) ;
    mux21_ni ix24924 (.Y (nx24923), .A0 (max_calc_comparator_first_inp1_7), .A1 (
             nx18064), .S0 (nx36285)) ;
    mux21_ni ix18065 (.Y (nx18064), .A0 (nx18060), .A1 (nx18028), .S0 (nx35973)
             ) ;
    mux21_ni ix18029 (.Y (nx18028), .A0 (max_calc_ans1_7), .A1 (
             label_1_output[7]), .S0 (nx35997)) ;
    mux21_ni ix24894 (.Y (nx24893), .A0 (nx13385), .A1 (max_calc_ans1_7), .S0 (
             nx35855)) ;
    mux21_ni ix18061 (.Y (nx18060), .A0 (max_calc_ans5_7), .A1 (max_calc_ans6_7)
             , .S0 (nx35997)) ;
    mux21_ni ix24904 (.Y (nx24903), .A0 (max_calc_ans6_7), .A1 (nx13385), .S0 (
             nx36025)) ;
    mux21_ni ix24914 (.Y (nx24913), .A0 (max_calc_ans5_7), .A1 (nx18050), .S0 (
             nx35751)) ;
    mux21 ix18051 (.Y (nx18050), .A0 (nx28040), .A1 (nx28044), .S0 (nx35863)) ;
    mux21_ni ix25034 (.Y (nx25033), .A0 (max_calc_comparator_first_inp2_6), .A1 (
             nx18224), .S0 (nx36285)) ;
    mux21_ni ix18225 (.Y (nx18224), .A0 (nx18220), .A1 (nx18132), .S0 (nx35973)
             ) ;
    mux21_ni ix18133 (.Y (nx18132), .A0 (max_calc_ans2_6), .A1 (
             label_2_output[6]), .S0 (nx35997)) ;
    mux21_ni ix24964 (.Y (nx24963), .A0 (nx18122), .A1 (max_calc_ans2_6), .S0 (
             nx35855)) ;
    mux21 ix18123 (.Y (nx18122), .A0 (nx33062), .A1 (nx33076), .S0 (nx35901)) ;
    mux21_ni ix18221 (.Y (nx18220), .A0 (max_calc_ans8_6), .A1 (max_calc_ans7_6)
             , .S0 (nx35997)) ;
    mux21_ni ix25024 (.Y (nx25023), .A0 (max_calc_ans7_6), .A1 (nx18122), .S0 (
             nx36025)) ;
    mux21_ni ix25014 (.Y (nx25013), .A0 (nx13386), .A1 (max_calc_ans8_6), .S0 (
             nx35871)) ;
    mux21_ni ix18201 (.Y (nx13386), .A0 (max_calc_comparator_first_inp2_6), .A1 (
             max_calc_comparator_first_inp1_6), .S0 (nx35907)) ;
    mux21_ni ix25004 (.Y (nx25003), .A0 (max_calc_comparator_first_inp1_6), .A1 (
             nx18186), .S0 (nx36285)) ;
    mux21_ni ix18187 (.Y (nx18186), .A0 (nx18182), .A1 (nx18150), .S0 (nx35973)
             ) ;
    mux21_ni ix18151 (.Y (nx18150), .A0 (max_calc_ans1_6), .A1 (
             label_1_output[6]), .S0 (nx35997)) ;
    mux21_ni ix24974 (.Y (nx24973), .A0 (nx13386), .A1 (max_calc_ans1_6), .S0 (
             nx35855)) ;
    mux21_ni ix18183 (.Y (nx18182), .A0 (max_calc_ans5_6), .A1 (max_calc_ans6_6)
             , .S0 (nx35997)) ;
    mux21_ni ix24984 (.Y (nx24983), .A0 (max_calc_ans6_6), .A1 (nx13386), .S0 (
             nx36025)) ;
    mux21_ni ix24994 (.Y (nx24993), .A0 (max_calc_ans5_6), .A1 (nx18172), .S0 (
             nx35751)) ;
    mux21 ix18173 (.Y (nx18172), .A0 (nx28051), .A1 (nx28058), .S0 (nx35863)) ;
    xor2 ix18233 (.Y (nx18232), .A0 (nx33950), .A1 (
         max_calc_comparator_first_inp1_6)) ;
    xor2 ix33987 (.Y (nx33986), .A0 (max_calc_comparator_first_inp2_5), .A1 (
         max_calc_comparator_first_inp1_5)) ;
    mux21_ni ix25114 (.Y (nx25113), .A0 (max_calc_comparator_first_inp2_5), .A1 (
             nx18346), .S0 (nx36287)) ;
    mux21_ni ix18347 (.Y (nx18346), .A0 (nx18342), .A1 (nx18254), .S0 (nx35973)
             ) ;
    mux21_ni ix18255 (.Y (nx18254), .A0 (max_calc_ans2_5), .A1 (
             label_2_output[5]), .S0 (nx35997)) ;
    mux21_ni ix25044 (.Y (nx25043), .A0 (nx18244), .A1 (max_calc_ans2_5), .S0 (
             nx35855)) ;
    mux21 ix18245 (.Y (nx18244), .A0 (nx33093), .A1 (nx33104), .S0 (nx35901)) ;
    mux21_ni ix18343 (.Y (nx18342), .A0 (max_calc_ans8_5), .A1 (max_calc_ans7_5)
             , .S0 (nx35189)) ;
    mux21_ni ix25104 (.Y (nx25103), .A0 (max_calc_ans7_5), .A1 (nx18244), .S0 (
             nx36025)) ;
    mux21_ni ix25094 (.Y (nx25093), .A0 (nx13387), .A1 (max_calc_ans8_5), .S0 (
             nx35871)) ;
    mux21_ni ix18323 (.Y (nx13387), .A0 (max_calc_comparator_first_inp2_5), .A1 (
             max_calc_comparator_first_inp1_5), .S0 (nx35907)) ;
    mux21_ni ix25084 (.Y (nx25083), .A0 (max_calc_comparator_first_inp1_5), .A1 (
             nx18308), .S0 (nx36287)) ;
    mux21_ni ix18309 (.Y (nx18308), .A0 (nx18304), .A1 (nx18272), .S0 (nx35973)
             ) ;
    mux21_ni ix18273 (.Y (nx18272), .A0 (max_calc_ans1_5), .A1 (
             label_1_output[5]), .S0 (nx35189)) ;
    mux21_ni ix25054 (.Y (nx25053), .A0 (nx13387), .A1 (max_calc_ans1_5), .S0 (
             nx35857)) ;
    mux21_ni ix18305 (.Y (nx18304), .A0 (max_calc_ans5_5), .A1 (max_calc_ans6_5)
             , .S0 (nx35189)) ;
    mux21_ni ix25064 (.Y (nx25063), .A0 (max_calc_ans6_5), .A1 (nx13387), .S0 (
             nx36027)) ;
    mux21_ni ix25074 (.Y (nx25073), .A0 (max_calc_ans5_5), .A1 (nx18294), .S0 (
             nx35751)) ;
    mux21 ix18295 (.Y (nx18294), .A0 (nx28068), .A1 (nx28072), .S0 (nx35863)) ;
    mux21_ni ix25194 (.Y (nx25193), .A0 (max_calc_comparator_first_inp2_4), .A1 (
             nx18468), .S0 (nx36287)) ;
    mux21_ni ix18469 (.Y (nx18468), .A0 (nx18464), .A1 (nx18376), .S0 (nx35975)
             ) ;
    mux21_ni ix18377 (.Y (nx18376), .A0 (max_calc_ans2_4), .A1 (
             label_2_output[4]), .S0 (nx35189)) ;
    mux21_ni ix25124 (.Y (nx25123), .A0 (nx18366), .A1 (max_calc_ans2_4), .S0 (
             nx35857)) ;
    mux21 ix18367 (.Y (nx18366), .A0 (nx33118), .A1 (nx33132), .S0 (nx35901)) ;
    mux21_ni ix18465 (.Y (nx18464), .A0 (max_calc_ans8_4), .A1 (max_calc_ans7_4)
             , .S0 (nx35189)) ;
    mux21_ni ix25184 (.Y (nx25183), .A0 (max_calc_ans7_4), .A1 (nx18366), .S0 (
             nx36027)) ;
    mux21_ni ix25174 (.Y (nx25173), .A0 (nx13388), .A1 (max_calc_ans8_4), .S0 (
             nx35871)) ;
    mux21_ni ix18445 (.Y (nx13388), .A0 (max_calc_comparator_first_inp2_4), .A1 (
             max_calc_comparator_first_inp1_4), .S0 (nx35907)) ;
    mux21_ni ix25164 (.Y (nx25163), .A0 (max_calc_comparator_first_inp1_4), .A1 (
             nx18430), .S0 (nx36287)) ;
    mux21_ni ix18431 (.Y (nx18430), .A0 (nx18426), .A1 (nx18394), .S0 (nx35975)
             ) ;
    mux21_ni ix18395 (.Y (nx18394), .A0 (max_calc_ans1_4), .A1 (
             label_1_output[4]), .S0 (nx35189)) ;
    mux21_ni ix25134 (.Y (nx25133), .A0 (nx13388), .A1 (max_calc_ans1_4), .S0 (
             nx35857)) ;
    mux21_ni ix18427 (.Y (nx18426), .A0 (max_calc_ans5_4), .A1 (max_calc_ans6_4)
             , .S0 (nx35189)) ;
    mux21_ni ix25144 (.Y (nx25143), .A0 (max_calc_ans6_4), .A1 (nx13388), .S0 (
             nx36027)) ;
    mux21_ni ix25154 (.Y (nx25153), .A0 (max_calc_ans5_4), .A1 (nx18416), .S0 (
             nx35751)) ;
    mux21 ix18417 (.Y (nx18416), .A0 (nx28079), .A1 (nx28086), .S0 (nx35863)) ;
    xor2 ix18477 (.Y (nx18476), .A0 (nx34023), .A1 (
         max_calc_comparator_first_inp1_4)) ;
    xor2 ix34060 (.Y (nx34059), .A0 (max_calc_comparator_first_inp2_3), .A1 (
         max_calc_comparator_first_inp1_3)) ;
    mux21_ni ix25274 (.Y (nx25273), .A0 (max_calc_comparator_first_inp2_3), .A1 (
             nx18590), .S0 (nx36287)) ;
    mux21_ni ix18591 (.Y (nx18590), .A0 (nx18586), .A1 (nx18498), .S0 (nx35975)
             ) ;
    mux21_ni ix18499 (.Y (nx18498), .A0 (max_calc_ans2_3), .A1 (
             label_2_output[3]), .S0 (nx35999)) ;
    mux21_ni ix25204 (.Y (nx25203), .A0 (nx18488), .A1 (max_calc_ans2_3), .S0 (
             nx35857)) ;
    mux21 ix18489 (.Y (nx18488), .A0 (nx33149), .A1 (nx33160), .S0 (nx35901)) ;
    mux21_ni ix18587 (.Y (nx18586), .A0 (max_calc_ans8_3), .A1 (max_calc_ans7_3)
             , .S0 (nx35999)) ;
    mux21_ni ix25264 (.Y (nx25263), .A0 (max_calc_ans7_3), .A1 (nx18488), .S0 (
             nx36027)) ;
    mux21_ni ix25254 (.Y (nx25253), .A0 (nx13389), .A1 (max_calc_ans8_3), .S0 (
             nx35871)) ;
    mux21_ni ix18567 (.Y (nx13389), .A0 (max_calc_comparator_first_inp2_3), .A1 (
             max_calc_comparator_first_inp1_3), .S0 (nx35907)) ;
    mux21_ni ix25244 (.Y (nx25243), .A0 (max_calc_comparator_first_inp1_3), .A1 (
             nx18552), .S0 (nx36287)) ;
    mux21_ni ix18553 (.Y (nx18552), .A0 (nx18548), .A1 (nx18516), .S0 (nx35975)
             ) ;
    mux21_ni ix18517 (.Y (nx18516), .A0 (max_calc_ans1_3), .A1 (
             label_1_output[3]), .S0 (nx35999)) ;
    mux21_ni ix25214 (.Y (nx25213), .A0 (nx13389), .A1 (max_calc_ans1_3), .S0 (
             nx35857)) ;
    mux21_ni ix18549 (.Y (nx18548), .A0 (max_calc_ans5_3), .A1 (max_calc_ans6_3)
             , .S0 (nx35999)) ;
    mux21_ni ix25224 (.Y (nx25223), .A0 (max_calc_ans6_3), .A1 (nx13389), .S0 (
             nx36027)) ;
    mux21_ni ix25234 (.Y (nx25233), .A0 (max_calc_ans5_3), .A1 (nx18538), .S0 (
             nx35751)) ;
    mux21 ix18539 (.Y (nx18538), .A0 (nx28096), .A1 (nx28100), .S0 (nx35863)) ;
    mux21_ni ix25354 (.Y (nx25353), .A0 (max_calc_comparator_first_inp2_2), .A1 (
             nx18712), .S0 (nx36287)) ;
    mux21_ni ix18713 (.Y (nx18712), .A0 (nx18708), .A1 (nx18620), .S0 (nx35975)
             ) ;
    mux21_ni ix18621 (.Y (nx18620), .A0 (max_calc_ans2_2), .A1 (
             label_2_output[2]), .S0 (nx35999)) ;
    mux21_ni ix25284 (.Y (nx25283), .A0 (nx18610), .A1 (max_calc_ans2_2), .S0 (
             nx35857)) ;
    mux21 ix18611 (.Y (nx18610), .A0 (nx33174), .A1 (nx33188), .S0 (nx35901)) ;
    mux21_ni ix18709 (.Y (nx18708), .A0 (max_calc_ans8_2), .A1 (max_calc_ans7_2)
             , .S0 (nx35999)) ;
    mux21_ni ix25344 (.Y (nx25343), .A0 (max_calc_ans7_2), .A1 (nx18610), .S0 (
             nx36027)) ;
    mux21_ni ix25334 (.Y (nx25333), .A0 (nx13391), .A1 (max_calc_ans8_2), .S0 (
             nx35873)) ;
    mux21_ni ix18689 (.Y (nx13391), .A0 (max_calc_comparator_first_inp2_2), .A1 (
             max_calc_comparator_first_inp1_2), .S0 (nx35907)) ;
    mux21_ni ix25324 (.Y (nx25323), .A0 (max_calc_comparator_first_inp1_2), .A1 (
             nx18674), .S0 (nx36289)) ;
    mux21_ni ix18675 (.Y (nx18674), .A0 (nx18670), .A1 (nx18638), .S0 (nx35975)
             ) ;
    mux21_ni ix18639 (.Y (nx18638), .A0 (max_calc_ans1_2), .A1 (
             label_1_output[2]), .S0 (nx35999)) ;
    mux21_ni ix25294 (.Y (nx25293), .A0 (nx13391), .A1 (max_calc_ans1_2), .S0 (
             nx35857)) ;
    mux21_ni ix18671 (.Y (nx18670), .A0 (max_calc_ans5_2), .A1 (max_calc_ans6_2)
             , .S0 (nx36001)) ;
    mux21_ni ix25304 (.Y (nx25303), .A0 (max_calc_ans6_2), .A1 (nx13391), .S0 (
             nx36027)) ;
    mux21_ni ix25314 (.Y (nx25313), .A0 (max_calc_ans5_2), .A1 (nx18660), .S0 (
             nx35751)) ;
    mux21 ix18661 (.Y (nx18660), .A0 (nx28107), .A1 (nx28114), .S0 (nx35863)) ;
    xor2 ix18721 (.Y (nx18720), .A0 (nx34096), .A1 (
         max_calc_comparator_first_inp1_2)) ;
    mux21_ni ix25434 (.Y (nx25433), .A0 (max_calc_comparator_first_inp2_1), .A1 (
             nx18834), .S0 (nx36289)) ;
    mux21_ni ix18835 (.Y (nx18834), .A0 (nx18830), .A1 (nx18742), .S0 (nx35975)
             ) ;
    mux21_ni ix18743 (.Y (nx18742), .A0 (max_calc_ans2_1), .A1 (
             label_2_output[1]), .S0 (nx36001)) ;
    mux21_ni ix25364 (.Y (nx25363), .A0 (nx18732), .A1 (max_calc_ans2_1), .S0 (
             nx35859)) ;
    mux21 ix18733 (.Y (nx18732), .A0 (nx33203), .A1 (nx33214), .S0 (nx35903)) ;
    mux21_ni ix18831 (.Y (nx18830), .A0 (max_calc_ans8_1), .A1 (max_calc_ans7_1)
             , .S0 (nx36001)) ;
    mux21_ni ix25424 (.Y (nx25423), .A0 (max_calc_ans7_1), .A1 (nx18732), .S0 (
             nx36029)) ;
    mux21_ni ix25414 (.Y (nx25413), .A0 (nx13393), .A1 (max_calc_ans8_1), .S0 (
             nx35873)) ;
    mux21_ni ix18811 (.Y (nx13393), .A0 (max_calc_comparator_first_inp2_1), .A1 (
             max_calc_comparator_first_inp1_1), .S0 (nx35909)) ;
    mux21_ni ix25404 (.Y (nx25403), .A0 (max_calc_comparator_first_inp1_1), .A1 (
             nx18796), .S0 (nx36289)) ;
    mux21_ni ix18797 (.Y (nx18796), .A0 (nx18792), .A1 (nx18760), .S0 (nx35185)
             ) ;
    mux21_ni ix18761 (.Y (nx18760), .A0 (max_calc_ans1_1), .A1 (
             label_1_output[1]), .S0 (nx36001)) ;
    mux21_ni ix25374 (.Y (nx25373), .A0 (nx13393), .A1 (max_calc_ans1_1), .S0 (
             nx35859)) ;
    mux21_ni ix18793 (.Y (nx18792), .A0 (max_calc_ans5_1), .A1 (max_calc_ans6_1)
             , .S0 (nx36001)) ;
    mux21_ni ix25384 (.Y (nx25383), .A0 (max_calc_ans6_1), .A1 (nx13393), .S0 (
             nx36029)) ;
    mux21_ni ix25394 (.Y (nx25393), .A0 (max_calc_ans5_1), .A1 (nx18782), .S0 (
             nx35753)) ;
    mux21 ix18783 (.Y (nx18782), .A0 (nx28122), .A1 (nx28126), .S0 (nx35865)) ;
    xor2 ix18843 (.Y (nx18842), .A0 (max_calc_comparator_first_inp2_1), .A1 (
         nx34162)) ;
    mux21_ni ix25554 (.Y (nx25553), .A0 (max_calc_comparator_first_inp2_15), .A1 (
             nx19132), .S0 (nx36289)) ;
    mux21_ni ix19133 (.Y (nx19132), .A0 (nx19128), .A1 (nx19040), .S0 (nx35185)
             ) ;
    mux21_ni ix19041 (.Y (nx19040), .A0 (max_calc_ans2_15), .A1 (
             label_2_output[15]), .S0 (nx36001)) ;
    mux21_ni ix16664 (.Y (nx16663), .A0 (label_2_output[15]), .A1 (
             label_2_input_15), .S0 (nx35609)) ;
    mux21_ni ix4889 (.Y (nx4888), .A0 (nx4884), .A1 (
             label_2_input_state_machine_15), .S0 (nx35171)) ;
    mux21_ni ix15824 (.Y (nx15823), .A0 (label_2_input_state_machine_15), .A1 (
             mdr_data_out[31]), .S0 (nx35601)) ;
    xor2 ix34183 (.Y (nx34182), .A0 (nx28594), .A1 (label_2_output[15])) ;
    mux21_ni ix25484 (.Y (nx25483), .A0 (nx19030), .A1 (max_calc_ans2_15), .S0 (
             nx35859)) ;
    mux21 ix19031 (.Y (nx19030), .A0 (nx33232), .A1 (nx33257), .S0 (nx35903)) ;
    mux21_ni ix19129 (.Y (nx19128), .A0 (max_calc_ans8_15), .A1 (
             max_calc_ans7_15), .S0 (nx36001)) ;
    mux21_ni ix25544 (.Y (nx25543), .A0 (max_calc_ans7_15), .A1 (nx19030), .S0 (
             nx36029)) ;
    mux21_ni ix25534 (.Y (nx25533), .A0 (nx13395), .A1 (max_calc_ans8_15), .S0 (
             nx35873)) ;
    mux21_ni ix19109 (.Y (nx13395), .A0 (max_calc_comparator_first_inp2_15), .A1 (
             max_calc_comparator_first_inp1_15), .S0 (nx35909)) ;
    mux21_ni ix25524 (.Y (nx25523), .A0 (max_calc_comparator_first_inp1_15), .A1 (
             nx19094), .S0 (nx36289)) ;
    mux21_ni ix19095 (.Y (nx19094), .A0 (nx19090), .A1 (nx19058), .S0 (nx35185)
             ) ;
    mux21_ni ix19059 (.Y (nx19058), .A0 (max_calc_ans1_15), .A1 (
             label_1_output[15]), .S0 (nx35191)) ;
    mux21_ni ix17514 (.Y (nx17513), .A0 (label_1_output[15]), .A1 (
             label_1_input_15), .S0 (nx35609)) ;
    mux21_ni ix6227 (.Y (nx6226), .A0 (nx6222), .A1 (
             label_1_input_state_machine_15), .S0 (nx35171)) ;
    mux21_ni ix16674 (.Y (nx16673), .A0 (label_1_input_state_machine_15), .A1 (
             mdr_data_out[15]), .S0 (nx35601)) ;
    xor2 ix34210 (.Y (nx34209), .A0 (nx26634), .A1 (label_1_output[15])) ;
    mux21_ni ix25494 (.Y (nx25493), .A0 (nx13395), .A1 (max_calc_ans1_15), .S0 (
             nx35859)) ;
    mux21_ni ix19091 (.Y (nx19090), .A0 (max_calc_ans5_15), .A1 (
             max_calc_ans6_15), .S0 (nx35191)) ;
    mux21_ni ix25504 (.Y (nx25503), .A0 (max_calc_ans6_15), .A1 (nx13395), .S0 (
             nx36029)) ;
    mux21_ni ix25514 (.Y (nx25513), .A0 (max_calc_ans5_15), .A1 (nx19080), .S0 (
             nx35753)) ;
    mux21 ix19081 (.Y (nx19080), .A0 (nx28137), .A1 (nx28155), .S0 (nx35865)) ;
    nor04 ix34227 (.Y (nx6342), .A0 (nx35737), .A1 (nx26180), .A2 (nx26203), .A3 (
          nx35711)) ;
    nand02 ix6341 (.Y (nx35711), .A0 (nx35191), .A1 (nx26188)) ;
    mux21_ni ix25574 (.Y (nx25573), .A0 (answer[1]), .A1 (nx13393), .S0 (nx35741
             )) ;
    mux21_ni ix25584 (.Y (nx25583), .A0 (answer[2]), .A1 (nx13391), .S0 (nx35741
             )) ;
    mux21_ni ix25594 (.Y (nx25593), .A0 (answer[3]), .A1 (nx13389), .S0 (nx35741
             )) ;
    mux21_ni ix25604 (.Y (nx25603), .A0 (answer[4]), .A1 (nx13388), .S0 (nx35741
             )) ;
    mux21_ni ix25614 (.Y (nx25613), .A0 (answer[5]), .A1 (nx13387), .S0 (nx35741
             )) ;
    mux21_ni ix25624 (.Y (nx25623), .A0 (answer[6]), .A1 (nx13386), .S0 (nx35743
             )) ;
    mux21_ni ix25634 (.Y (nx25633), .A0 (answer[7]), .A1 (nx13385), .S0 (nx35743
             )) ;
    mux21_ni ix25644 (.Y (nx25643), .A0 (answer[8]), .A1 (nx13383), .S0 (nx35743
             )) ;
    mux21_ni ix25654 (.Y (nx25653), .A0 (answer[9]), .A1 (nx13381), .S0 (nx35743
             )) ;
    mux21_ni ix25664 (.Y (nx25663), .A0 (answer[10]), .A1 (nx13379), .S0 (
             nx35743)) ;
    mux21_ni ix25674 (.Y (nx25673), .A0 (answer[11]), .A1 (nx13377), .S0 (
             nx35743)) ;
    mux21_ni ix25684 (.Y (nx25683), .A0 (answer[12]), .A1 (nx13376), .S0 (
             nx35743)) ;
    mux21_ni ix25694 (.Y (nx25693), .A0 (answer[13]), .A1 (nx13375), .S0 (
             nx35745)) ;
    mux21_ni ix25704 (.Y (nx25703), .A0 (answer[14]), .A1 (nx13371), .S0 (
             nx35745)) ;
    mux21_ni ix25714 (.Y (nx25713), .A0 (answer[15]), .A1 (nx13395), .S0 (
             nx35745)) ;
    and02 ix191 (.Y (nx190), .A0 (nx12893), .A1 (nx25907)) ;
    nor02ii ix19277 (.Y (nx19276), .A0 (nx38), .A1 (nx12887)) ;
    nor02ii ix19241 (.Y (nx19240), .A0 (nx34380), .A1 (nx26129)) ;
    nor02ii ix34381 (.Y (nx34380), .A0 (nx19232), .A1 (nx12879)) ;
    and02 ix34584 (.Y (nx34585), .A0 (nx30681), .A1 (nx35721)) ;
    and02 ix34586 (.Y (nx34587), .A0 (nx30681), .A1 (nx35721)) ;
    and02 ix34616 (.Y (nx34617), .A0 (nx28752), .A1 (nx35725)) ;
    and02 ix34618 (.Y (nx34619), .A0 (nx28752), .A1 (nx35725)) ;
    and02 ix34648 (.Y (nx34649), .A0 (nx28309), .A1 (nx35729)) ;
    and02 ix34650 (.Y (nx34651), .A0 (nx28309), .A1 (nx35729)) ;
    and02 ix34680 (.Y (nx34681), .A0 (nx26349), .A1 (nx35733)) ;
    and02 ix34682 (.Y (nx34683), .A0 (nx26349), .A1 (nx35733)) ;
    and02 ix34860 (.Y (nx34861), .A0 (nx26828), .A1 (nx35757)) ;
    and02 ix34862 (.Y (nx34863), .A0 (nx26828), .A1 (nx35757)) ;
    and02 ix34892 (.Y (nx34893), .A0 (nx27267), .A1 (nx35761)) ;
    and02 ix34894 (.Y (nx34895), .A0 (nx27267), .A1 (nx35761)) ;
    and02 ix34952 (.Y (nx34953), .A0 (nx29195), .A1 (nx35765)) ;
    and02 ix34954 (.Y (nx34955), .A0 (nx29195), .A1 (nx35765)) ;
    and02 ix34984 (.Y (nx34985), .A0 (nx29636), .A1 (nx35769)) ;
    and02 ix34986 (.Y (nx34987), .A0 (nx29636), .A1 (nx35769)) ;
    and02 ix35024 (.Y (nx35025), .A0 (nx31124), .A1 (nx35773)) ;
    and02 ix35026 (.Y (nx35027), .A0 (nx31124), .A1 (nx35773)) ;
    and02 ix35056 (.Y (nx35057), .A0 (nx31563), .A1 (nx35777)) ;
    and02 ix35058 (.Y (nx35059), .A0 (nx31563), .A1 (nx35777)) ;
    inv02 ix35712 (.Y (nx35713), .A (nx35149)) ;
    inv02 ix35714 (.Y (nx35715), .A (nx35149)) ;
    inv02 ix35716 (.Y (nx35717), .A (nx35149)) ;
    inv01 ix35718 (.Y (nx35719), .A (nx30685)) ;
    inv01 ix35720 (.Y (nx35721), .A (nx30685)) ;
    inv01 ix35722 (.Y (nx35723), .A (nx28756)) ;
    inv01 ix35724 (.Y (nx35725), .A (nx28756)) ;
    inv01 ix35726 (.Y (nx35727), .A (nx28313)) ;
    inv01 ix35728 (.Y (nx35729), .A (nx28313)) ;
    inv01 ix35730 (.Y (nx35731), .A (nx26353)) ;
    inv01 ix35732 (.Y (nx35733), .A (nx26353)) ;
    inv02 ix35734 (.Y (nx35735), .A (nx36389)) ;
    inv02 ix35736 (.Y (nx35737), .A (nx36389)) ;
    inv01 ix35738 (.Y (nx35739), .A (nx6342)) ;
    inv02 ix35740 (.Y (nx35741), .A (nx35739)) ;
    inv02 ix35742 (.Y (nx35743), .A (nx35739)) ;
    inv02 ix35744 (.Y (nx35745), .A (nx35739)) ;
    inv02 ix35746 (.Y (nx35747), .A (nx26675)) ;
    inv02 ix35748 (.Y (nx35749), .A (nx36381)) ;
    inv02 ix35750 (.Y (nx35751), .A (nx36381)) ;
    inv02 ix35752 (.Y (nx35753), .A (nx36381)) ;
    inv01 ix35754 (.Y (nx35755), .A (nx26832)) ;
    inv01 ix35756 (.Y (nx35757), .A (nx26832)) ;
    inv01 ix35758 (.Y (nx35759), .A (nx27271)) ;
    inv01 ix35760 (.Y (nx35761), .A (nx27271)) ;
    inv01 ix35762 (.Y (nx35763), .A (nx29199)) ;
    inv01 ix35764 (.Y (nx35765), .A (nx29199)) ;
    inv01 ix35766 (.Y (nx35767), .A (nx29640)) ;
    inv01 ix35768 (.Y (nx35769), .A (nx29640)) ;
    inv01 ix35770 (.Y (nx35771), .A (nx31128)) ;
    inv01 ix35772 (.Y (nx35773), .A (nx31128)) ;
    inv01 ix35774 (.Y (nx35775), .A (nx31567)) ;
    inv01 ix35776 (.Y (nx35777), .A (nx31567)) ;
    inv02 ix35778 (.Y (nx35779), .A (state[1])) ;
    inv02 ix35780 (.Y (nx35781), .A (state[1])) ;
    inv02 ix35782 (.Y (nx35783), .A (state[2])) ;
    inv02 ix35784 (.Y (nx35785), .A (state[2])) ;
    buf02 ix35786 (.Y (nx35787), .A (nx25874)) ;
    buf02 ix35788 (.Y (nx35789), .A (nx25874)) ;
    inv01 ix35790 (.Y (nx35791), .A (sub_state[2])) ;
    inv01 ix35792 (.Y (nx35793), .A (sub_state[2])) ;
    buf02 ix35794 (.Y (nx35795), .A (nx25949)) ;
    buf02 ix35796 (.Y (nx35797), .A (nx25949)) ;
    inv02 ix35798 (.Y (nx35799), .A (nx34499)) ;
    inv02 ix35800 (.Y (nx35801), .A (nx34499)) ;
    buf02 ix35802 (.Y (nx35803), .A (nx26323)) ;
    buf02 ix35804 (.Y (nx35805), .A (nx26323)) ;
    buf02 ix35806 (.Y (nx35807), .A (nx26802)) ;
    buf02 ix35808 (.Y (nx35809), .A (nx26802)) ;
    buf02 ix35810 (.Y (nx35811), .A (nx27241)) ;
    buf02 ix35812 (.Y (nx35813), .A (nx27241)) ;
    buf02 ix35814 (.Y (nx35815), .A (nx28283)) ;
    buf02 ix35816 (.Y (nx35817), .A (nx28283)) ;
    buf02 ix35818 (.Y (nx35819), .A (nx28726)) ;
    buf02 ix35820 (.Y (nx35821), .A (nx28726)) ;
    buf02 ix35822 (.Y (nx35823), .A (nx29169)) ;
    buf02 ix35824 (.Y (nx35825), .A (nx29169)) ;
    buf02 ix35826 (.Y (nx35827), .A (nx29610)) ;
    buf02 ix35828 (.Y (nx35829), .A (nx29610)) ;
    buf02 ix35830 (.Y (nx35831), .A (nx30655)) ;
    buf02 ix35832 (.Y (nx35833), .A (nx30655)) ;
    buf02 ix35834 (.Y (nx35835), .A (nx31098)) ;
    buf02 ix35836 (.Y (nx35837), .A (nx31098)) ;
    buf02 ix35838 (.Y (nx35839), .A (nx31537)) ;
    buf02 ix35840 (.Y (nx35841), .A (nx31537)) ;
    inv02 ix35842 (.Y (nx35843), .A (nx34737)) ;
    inv02 ix35844 (.Y (nx35845), .A (nx34737)) ;
    inv02 ix35846 (.Y (nx35847), .A (nx34737)) ;
    inv01 ix35848 (.Y (nx35849), .A (nx34821)) ;
    inv02 ix35850 (.Y (nx35851), .A (nx35849)) ;
    inv02 ix35852 (.Y (nx35853), .A (nx35849)) ;
    inv02 ix35854 (.Y (nx35855), .A (nx35849)) ;
    inv02 ix35856 (.Y (nx35857), .A (nx35849)) ;
    inv02 ix35858 (.Y (nx35859), .A (nx35849)) ;
    inv02 ix35860 (.Y (nx35861), .A (nx9490)) ;
    inv02 ix35862 (.Y (nx35863), .A (nx9490)) ;
    inv02 ix35864 (.Y (nx35865), .A (nx9490)) ;
    inv01 ix35866 (.Y (nx35867), .A (nx34905)) ;
    inv02 ix35868 (.Y (nx35869), .A (nx35867)) ;
    inv02 ix35870 (.Y (nx35871), .A (nx35867)) ;
    inv02 ix35872 (.Y (nx35873), .A (nx35867)) ;
    inv01 ix35874 (.Y (nx35875), .A (nx34913)) ;
    inv02 ix35876 (.Y (nx35877), .A (nx35875)) ;
    inv02 ix35878 (.Y (nx35879), .A (nx35875)) ;
    inv02 ix35880 (.Y (nx35881), .A (nx35875)) ;
    inv02 ix35882 (.Y (nx35883), .A (nx35875)) ;
    inv02 ix35884 (.Y (nx35885), .A (nx35875)) ;
    inv02 ix35886 (.Y (nx35887), .A (nx12690)) ;
    inv02 ix35888 (.Y (nx35889), .A (nx12690)) ;
    inv02 ix35890 (.Y (nx35891), .A (nx12690)) ;
    inv02 ix35892 (.Y (nx35893), .A (nx15874)) ;
    inv02 ix35894 (.Y (nx35895), .A (nx15874)) ;
    inv02 ix35896 (.Y (nx35897), .A (nx15874)) ;
    inv02 ix35898 (.Y (nx35899), .A (nx17138)) ;
    inv02 ix35900 (.Y (nx35901), .A (nx17138)) ;
    inv02 ix35902 (.Y (nx35903), .A (nx17138)) ;
    inv02 ix35904 (.Y (nx35905), .A (nx13373)) ;
    inv02 ix35906 (.Y (nx35907), .A (nx13373)) ;
    inv02 ix35908 (.Y (nx35909), .A (nx13373)) ;
    inv02 ix35910 (.Y (nx35911), .A (done)) ;
    inv02 ix35912 (.Y (nx35913), .A (done)) ;
    inv02 ix35914 (.Y (nx35915), .A (done)) ;
    inv02 ix35916 (.Y (nx35917), .A (done)) ;
    inv02 ix35918 (.Y (nx35919), .A (nx36307)) ;
    inv02 ix35920 (.Y (nx35921), .A (nx36307)) ;
    inv02 ix35922 (.Y (nx35923), .A (nx36307)) ;
    inv02 ix35924 (.Y (nx35925), .A (nx36309)) ;
    inv02 ix35926 (.Y (nx35927), .A (nx36309)) ;
    inv02 ix35928 (.Y (nx35929), .A (nx36309)) ;
    inv02 ix35930 (.Y (nx35931), .A (nx36309)) ;
    inv02 ix35932 (.Y (nx35933), .A (nx36309)) ;
    inv02 ix35934 (.Y (nx35935), .A (nx36309)) ;
    inv02 ix35936 (.Y (nx35937), .A (nx36309)) ;
    inv02 ix35938 (.Y (nx35939), .A (nx36311)) ;
    inv02 ix35940 (.Y (nx35941), .A (nx36311)) ;
    inv02 ix35942 (.Y (nx35943), .A (nx36311)) ;
    inv02 ix35944 (.Y (nx35945), .A (nx36311)) ;
    inv02 ix35946 (.Y (nx35947), .A (nx36311)) ;
    inv02 ix35948 (.Y (nx35949), .A (nx36311)) ;
    inv02 ix35950 (.Y (nx35951), .A (nx36311)) ;
    inv02 ix35952 (.Y (nx35953), .A (nx36313)) ;
    inv02 ix35954 (.Y (nx35955), .A (nx36313)) ;
    inv02 ix35956 (.Y (nx35957), .A (nx36313)) ;
    inv02 ix35958 (.Y (nx35959), .A (nx36301)) ;
    inv02 ix35960 (.Y (nx35961), .A (nx36301)) ;
    inv02 ix35962 (.Y (nx35963), .A (nx36301)) ;
    inv02 ix35964 (.Y (nx35965), .A (nx36301)) ;
    inv02 ix35966 (.Y (nx35967), .A (nx36301)) ;
    inv02 ix35968 (.Y (nx35969), .A (nx36301)) ;
    inv02 ix35970 (.Y (nx35971), .A (nx36301)) ;
    inv02 ix35972 (.Y (nx35973), .A (nx35735)) ;
    inv02 ix35974 (.Y (nx35975), .A (nx35735)) ;
    inv02 ix35976 (.Y (nx35977), .A (nx36331)) ;
    inv02 ix35978 (.Y (nx35979), .A (nx36331)) ;
    inv02 ix35980 (.Y (nx35981), .A (nx36331)) ;
    inv02 ix35982 (.Y (nx35983), .A (nx36331)) ;
    inv02 ix35984 (.Y (nx35985), .A (nx36333)) ;
    inv02 ix35986 (.Y (nx35987), .A (nx36333)) ;
    inv02 ix35988 (.Y (nx35989), .A (nx36333)) ;
    inv02 ix35990 (.Y (nx35991), .A (nx36333)) ;
    inv02 ix35992 (.Y (nx35993), .A (nx36333)) ;
    inv02 ix35994 (.Y (nx35995), .A (nx36333)) ;
    inv02 ix35996 (.Y (nx35997), .A (nx36333)) ;
    inv02 ix35998 (.Y (nx35999), .A (nx36335)) ;
    inv02 ix36000 (.Y (nx36001), .A (nx36335)) ;
    inv02 ix36002 (.Y (nx36003), .A (nx36327)) ;
    inv02 ix36004 (.Y (nx36005), .A (nx36327)) ;
    inv02 ix36006 (.Y (nx36007), .A (nx36329)) ;
    inv02 ix36008 (.Y (nx36009), .A (nx36329)) ;
    inv02 ix36010 (.Y (nx36011), .A (
          booth_booth_integrtaion_0_shift_reg_output_0)) ;
    inv02 ix36012 (.Y (nx36013), .A (
          booth_booth_integrtaion_0_shift_reg_output_0)) ;
    inv02 ix36014 (.Y (nx36015), .A (
          booth_booth_integrtaion_0_shift_reg_output_0)) ;
    inv02 ix36016 (.Y (nx36017), .A (
          booth_booth_integrtaion_0_shift_reg_output_0)) ;
    inv01 ix36018 (.Y (nx36019), .A (nx35289)) ;
    inv02 ix36020 (.Y (nx36021), .A (nx36019)) ;
    inv02 ix36022 (.Y (nx36023), .A (nx36019)) ;
    inv02 ix36024 (.Y (nx36025), .A (nx36019)) ;
    inv02 ix36026 (.Y (nx36027), .A (nx36019)) ;
    inv02 ix36028 (.Y (nx36029), .A (nx36019)) ;
    inv02 ix36030 (.Y (nx36031), .A (nx36341)) ;
    inv02 ix36032 (.Y (nx36033), .A (nx36341)) ;
    inv02 ix36034 (.Y (nx36035), .A (nx36343)) ;
    inv02 ix36036 (.Y (nx36037), .A (nx36343)) ;
    inv02 ix36038 (.Y (nx36039), .A (
          booth_booth_integrtaion_8_shift_reg_output_0)) ;
    inv02 ix36040 (.Y (nx36041), .A (
          booth_booth_integrtaion_8_shift_reg_output_0)) ;
    inv02 ix36042 (.Y (nx36043), .A (
          booth_booth_integrtaion_8_shift_reg_output_0)) ;
    inv02 ix36044 (.Y (nx36045), .A (
          booth_booth_integrtaion_8_shift_reg_output_0)) ;
    inv02 ix36046 (.Y (nx36047), .A (nx36345)) ;
    inv02 ix36048 (.Y (nx36049), .A (nx36345)) ;
    inv02 ix36050 (.Y (nx36051), .A (nx36347)) ;
    inv02 ix36052 (.Y (nx36053), .A (nx36347)) ;
    inv02 ix36054 (.Y (nx36055), .A (
          booth_booth_integrtaion_9_shift_reg_output_0)) ;
    inv02 ix36056 (.Y (nx36057), .A (
          booth_booth_integrtaion_9_shift_reg_output_0)) ;
    inv02 ix36058 (.Y (nx36059), .A (
          booth_booth_integrtaion_9_shift_reg_output_0)) ;
    inv02 ix36060 (.Y (nx36061), .A (
          booth_booth_integrtaion_9_shift_reg_output_0)) ;
    inv02 ix36062 (.Y (nx36063), .A (nx36337)) ;
    inv02 ix36064 (.Y (nx36065), .A (nx36337)) ;
    inv02 ix36066 (.Y (nx36067), .A (nx36339)) ;
    inv02 ix36068 (.Y (nx36069), .A (nx36339)) ;
    inv02 ix36070 (.Y (nx36071), .A (nx36339)) ;
    inv02 ix36072 (.Y (nx36073), .A (nx36339)) ;
    inv02 ix36074 (.Y (nx36075), .A (nx36339)) ;
    inv02 ix36076 (.Y (nx36077), .A (nx36323)) ;
    inv02 ix36078 (.Y (nx36079), .A (nx36323)) ;
    inv02 ix36080 (.Y (nx36081), .A (nx36325)) ;
    inv02 ix36082 (.Y (nx36083), .A (nx36325)) ;
    inv02 ix36084 (.Y (nx36085), .A (
          booth_booth_integrtaion_1_shift_reg_output_0)) ;
    inv02 ix36086 (.Y (nx36087), .A (
          booth_booth_integrtaion_1_shift_reg_output_0)) ;
    inv02 ix36088 (.Y (nx36089), .A (
          booth_booth_integrtaion_1_shift_reg_output_0)) ;
    inv02 ix36090 (.Y (nx36091), .A (
          booth_booth_integrtaion_1_shift_reg_output_0)) ;
    inv02 ix36092 (.Y (nx36093), .A (nx36319)) ;
    inv02 ix36094 (.Y (nx36095), .A (nx36319)) ;
    inv02 ix36096 (.Y (nx36097), .A (nx36321)) ;
    inv02 ix36098 (.Y (nx36099), .A (nx36321)) ;
    inv02 ix36100 (.Y (nx36101), .A (
          booth_booth_integrtaion_2_shift_reg_output_0)) ;
    inv02 ix36102 (.Y (nx36103), .A (
          booth_booth_integrtaion_2_shift_reg_output_0)) ;
    inv02 ix36104 (.Y (nx36105), .A (
          booth_booth_integrtaion_2_shift_reg_output_0)) ;
    inv02 ix36106 (.Y (nx36107), .A (
          booth_booth_integrtaion_2_shift_reg_output_0)) ;
    inv02 ix36108 (.Y (nx36109), .A (nx36349)) ;
    inv02 ix36110 (.Y (nx36111), .A (nx36349)) ;
    inv02 ix36112 (.Y (nx36113), .A (nx36351)) ;
    inv02 ix36114 (.Y (nx36115), .A (nx36351)) ;
    inv02 ix36116 (.Y (nx36117), .A (
          booth_booth_integrtaion_4_shift_reg_output_0)) ;
    inv02 ix36118 (.Y (nx36119), .A (
          booth_booth_integrtaion_4_shift_reg_output_0)) ;
    inv02 ix36120 (.Y (nx36121), .A (
          booth_booth_integrtaion_4_shift_reg_output_0)) ;
    inv02 ix36122 (.Y (nx36123), .A (
          booth_booth_integrtaion_4_shift_reg_output_0)) ;
    inv02 ix36124 (.Y (nx36125), .A (nx29498)) ;
    inv02 ix36126 (.Y (nx36127), .A (nx29498)) ;
    inv02 ix36128 (.Y (nx36129), .A (nx29498)) ;
    inv02 ix36130 (.Y (nx36131), .A (nx36353)) ;
    inv02 ix36132 (.Y (nx36133), .A (nx36353)) ;
    inv02 ix36134 (.Y (nx36135), .A (nx36355)) ;
    inv02 ix36136 (.Y (nx36137), .A (nx36355)) ;
    inv02 ix36138 (.Y (nx36139), .A (
          booth_booth_integrtaion_5_shift_reg_output_0)) ;
    inv02 ix36140 (.Y (nx36141), .A (
          booth_booth_integrtaion_5_shift_reg_output_0)) ;
    inv02 ix36142 (.Y (nx36143), .A (
          booth_booth_integrtaion_5_shift_reg_output_0)) ;
    inv02 ix36144 (.Y (nx36145), .A (
          booth_booth_integrtaion_5_shift_reg_output_0)) ;
    inv02 ix36146 (.Y (nx36147), .A (nx36315)) ;
    inv02 ix36148 (.Y (nx36149), .A (nx36315)) ;
    inv02 ix36150 (.Y (nx36151), .A (nx36317)) ;
    inv02 ix36152 (.Y (nx36153), .A (nx36317)) ;
    inv02 ix36154 (.Y (nx36155), .A (
          booth_booth_integrtaion_3_shift_reg_output_0)) ;
    inv02 ix36156 (.Y (nx36157), .A (
          booth_booth_integrtaion_3_shift_reg_output_0)) ;
    inv02 ix36158 (.Y (nx36159), .A (
          booth_booth_integrtaion_3_shift_reg_output_0)) ;
    inv02 ix36160 (.Y (nx36161), .A (
          booth_booth_integrtaion_3_shift_reg_output_0)) ;
    inv02 ix36162 (.Y (nx36163), .A (nx36357)) ;
    inv02 ix36164 (.Y (nx36165), .A (nx36357)) ;
    inv02 ix36166 (.Y (nx36167), .A (nx36359)) ;
    inv02 ix36168 (.Y (nx36169), .A (nx36359)) ;
    inv02 ix36170 (.Y (nx36171), .A (
          booth_booth_integrtaion_6_shift_reg_output_0)) ;
    inv02 ix36172 (.Y (nx36173), .A (
          booth_booth_integrtaion_6_shift_reg_output_0)) ;
    inv02 ix36174 (.Y (nx36175), .A (
          booth_booth_integrtaion_6_shift_reg_output_0)) ;
    inv02 ix36176 (.Y (nx36177), .A (
          booth_booth_integrtaion_6_shift_reg_output_0)) ;
    inv02 ix36178 (.Y (nx36179), .A (nx36361)) ;
    inv02 ix36180 (.Y (nx36181), .A (nx36361)) ;
    inv02 ix36182 (.Y (nx36183), .A (nx36363)) ;
    inv02 ix36184 (.Y (nx36185), .A (nx36363)) ;
    inv02 ix36186 (.Y (nx36187), .A (
          booth_booth_integrtaion_7_shift_reg_output_0)) ;
    inv02 ix36188 (.Y (nx36189), .A (
          booth_booth_integrtaion_7_shift_reg_output_0)) ;
    inv02 ix36190 (.Y (nx36191), .A (
          booth_booth_integrtaion_7_shift_reg_output_0)) ;
    inv02 ix36192 (.Y (nx36193), .A (
          booth_booth_integrtaion_7_shift_reg_output_0)) ;
    inv02 ix36194 (.Y (nx36195), .A (nx29498)) ;
    inv02 ix36196 (.Y (nx36197), .A (nx29498)) ;
    inv02 ix36198 (.Y (nx36199), .A (nx29498)) ;
    inv02 ix36200 (.Y (nx36201), .A (nx36365)) ;
    inv02 ix36202 (.Y (nx36203), .A (nx36365)) ;
    inv02 ix36204 (.Y (nx36205), .A (nx36365)) ;
    inv02 ix36206 (.Y (nx36207), .A (nx36365)) ;
    inv02 ix36208 (.Y (nx36209), .A (nx36367)) ;
    inv02 ix36210 (.Y (nx36211), .A (nx36367)) ;
    inv02 ix36212 (.Y (nx36213), .A (nx36367)) ;
    inv02 ix36214 (.Y (nx36215), .A (nx36367)) ;
    inv02 ix36216 (.Y (nx36217), .A (nx36367)) ;
    inv02 ix36218 (.Y (nx36219), .A (nx36367)) ;
    inv02 ix36220 (.Y (nx36221), .A (nx36367)) ;
    inv02 ix36222 (.Y (nx36223), .A (nx36369)) ;
    inv02 ix36224 (.Y (nx36225), .A (nx36369)) ;
    inv02 ix36226 (.Y (nx36227), .A (nx36369)) ;
    inv02 ix36228 (.Y (nx36229), .A (nx36369)) ;
    inv02 ix36230 (.Y (nx36231), .A (nx36369)) ;
    inv02 ix36232 (.Y (nx36233), .A (nx36369)) ;
    inv02 ix36234 (.Y (nx36235), .A (nx36369)) ;
    inv02 ix36236 (.Y (nx36237), .A (nx36371)) ;
    inv02 ix36238 (.Y (nx36239), .A (nx36371)) ;
    inv02 ix36240 (.Y (nx36241), .A (nx36373)) ;
    inv02 ix36242 (.Y (nx36243), .A (nx36373)) ;
    inv02 ix36244 (.Y (nx36245), .A (nx36373)) ;
    inv02 ix36246 (.Y (nx36247), .A (nx36373)) ;
    inv02 ix36248 (.Y (nx36249), .A (nx36375)) ;
    inv02 ix36250 (.Y (nx36251), .A (nx36375)) ;
    inv02 ix36252 (.Y (nx36253), .A (nx36375)) ;
    inv02 ix36254 (.Y (nx36255), .A (nx36375)) ;
    inv02 ix36256 (.Y (nx36257), .A (nx36375)) ;
    inv02 ix36258 (.Y (nx36259), .A (nx36375)) ;
    inv02 ix36260 (.Y (nx36261), .A (nx36375)) ;
    inv02 ix36262 (.Y (nx36263), .A (nx36377)) ;
    inv02 ix36264 (.Y (nx36265), .A (nx36377)) ;
    inv02 ix36266 (.Y (nx36267), .A (nx36377)) ;
    inv02 ix36268 (.Y (nx36269), .A (nx36377)) ;
    inv02 ix36270 (.Y (nx36271), .A (nx36377)) ;
    inv02 ix36272 (.Y (nx36273), .A (nx36377)) ;
    inv02 ix36274 (.Y (nx36275), .A (nx36377)) ;
    inv02 ix36276 (.Y (nx36277), .A (nx36379)) ;
    inv02 ix36278 (.Y (nx36279), .A (nx36379)) ;
    inv02 ix36280 (.Y (nx36281), .A (nx36385)) ;
    inv02 ix36282 (.Y (nx36283), .A (nx36385)) ;
    inv02 ix36284 (.Y (nx36285), .A (nx36385)) ;
    inv02 ix36286 (.Y (nx36287), .A (nx36385)) ;
    inv02 ix36288 (.Y (nx36289), .A (nx36385)) ;
    inv02 ix36290 (.Y (nx36291), .A (nx36381)) ;
    inv02 ix36292 (.Y (nx36293), .A (nx36381)) ;
    inv02 ix36294 (.Y (nx36295), .A (nx36381)) ;
    inv02 ix36296 (.Y (nx36297), .A (nx36383)) ;
    inv02 ix36298 (.Y (nx36299), .A (nx35173)) ;
    inv02 ix36300 (.Y (nx36301), .A (nx35173)) ;
    inv02 ix36306 (.Y (nx36307), .A (nx35163)) ;
    inv02 ix36308 (.Y (nx36309), .A (nx35163)) ;
    inv02 ix36310 (.Y (nx36311), .A (nx35163)) ;
    inv02 ix36312 (.Y (nx36313), .A (nx35163)) ;
    inv02 ix36314 (.Y (nx36315), .A (nx35499)) ;
    inv02 ix36316 (.Y (nx36317), .A (nx35499)) ;
    inv02 ix36318 (.Y (nx36319), .A (nx35399)) ;
    inv02 ix36320 (.Y (nx36321), .A (nx35399)) ;
    inv02 ix36322 (.Y (nx36323), .A (nx35373)) ;
    inv02 ix36324 (.Y (nx36325), .A (nx35373)) ;
    inv02 ix36326 (.Y (nx36327), .A (nx35193)) ;
    inv02 ix36328 (.Y (nx36329), .A (nx35193)) ;
    inv02 ix36330 (.Y (nx36331), .A (nx35187)) ;
    inv02 ix36332 (.Y (nx36333), .A (nx35187)) ;
    inv02 ix36334 (.Y (nx36335), .A (nx35187)) ;
    inv02 ix36336 (.Y (nx36337), .A (nx36385)) ;
    inv02 ix36338 (.Y (nx36339), .A (nx36385)) ;
    inv02 ix36340 (.Y (nx36341), .A (nx35301)) ;
    inv02 ix36342 (.Y (nx36343), .A (nx35301)) ;
    inv02 ix36344 (.Y (nx36345), .A (nx35327)) ;
    inv02 ix36346 (.Y (nx36347), .A (nx35327)) ;
    inv02 ix36348 (.Y (nx36349), .A (nx35425)) ;
    inv02 ix36350 (.Y (nx36351), .A (nx35425)) ;
    inv02 ix36352 (.Y (nx36353), .A (nx35473)) ;
    inv02 ix36354 (.Y (nx36355), .A (nx35473)) ;
    inv02 ix36356 (.Y (nx36357), .A (nx35525)) ;
    inv02 ix36358 (.Y (nx36359), .A (nx35525)) ;
    inv02 ix36360 (.Y (nx36361), .A (nx35551)) ;
    inv02 ix36362 (.Y (nx36363), .A (nx35551)) ;
    inv02 ix36364 (.Y (nx36365), .A (nx35595)) ;
    inv02 ix36366 (.Y (nx36367), .A (nx35595)) ;
    inv02 ix36368 (.Y (nx36369), .A (nx35595)) ;
    inv02 ix36370 (.Y (nx36371), .A (nx35595)) ;
    inv02 ix36372 (.Y (nx36373), .A (nx35603)) ;
    inv02 ix36374 (.Y (nx36375), .A (nx35603)) ;
    inv02 ix36376 (.Y (nx36377), .A (nx35603)) ;
    inv02 ix36378 (.Y (nx36379), .A (nx35603)) ;
    inv02 ix36380 (.Y (nx36381), .A (nx35747)) ;
    inv02 ix36382 (.Y (nx36383), .A (nx35747)) ;
    inv02 ix36384 (.Y (nx36385), .A (nx6352)) ;
    inv02 ix36386 (.Y (nx36387), .A (enable_decoder_dst_booth)) ;
    inv02 ix36388 (.Y (nx36389), .A (max_calc_state_2)) ;
    inv02 ix36390 (.Y (nx36391), .A (nx26669)) ;
    inv02 ix36392 (.Y (nx36393), .A (nx26675)) ;
endmodule

